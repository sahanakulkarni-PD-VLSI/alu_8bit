VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu_8bit
  CLASS BLOCK ;
  FOREIGN alu_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.820 BY 65.540 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.480 10.640 15.080 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.405 10.640 26.005 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.330 10.640 36.930 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.255 10.640 47.855 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.815 49.460 20.415 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.690 49.460 31.290 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.565 49.460 42.165 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 51.440 49.460 53.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.180 10.640 11.780 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.105 10.640 22.705 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.030 10.640 33.630 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.955 10.640 44.555 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.515 49.460 17.115 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.390 49.460 27.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 37.265 49.460 38.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 48.140 49.460 49.740 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 50.820 23.840 54.820 24.440 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 61.540 39.010 65.540 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 61.540 32.570 65.540 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 61.540 19.690 65.540 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 50.820 20.440 54.820 21.040 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 50.820 27.240 54.820 27.840 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 61.540 42.230 65.540 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 61.540 29.350 65.540 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END b[7]
  PIN cin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END cin
  PIN cout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END cout
  PIN op[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END op[0]
  PIN op[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 50.820 34.040 54.820 34.640 ;
    END
  END op[1]
  PIN op[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 50.820 40.840 54.820 41.440 ;
    END
  END op[2]
  PIN result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END result[0]
  PIN result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 50.820 30.640 54.820 31.240 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 50.820 37.440 54.820 38.040 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 61.540 26.130 65.540 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END result[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 49.410 54.485 ;
      LAYER li1 ;
        RECT 5.520 10.795 49.220 54.485 ;
      LAYER met1 ;
        RECT 4.210 10.640 49.220 54.640 ;
      LAYER met2 ;
        RECT 4.230 61.260 19.130 61.540 ;
        RECT 19.970 61.260 25.570 61.540 ;
        RECT 26.410 61.260 28.790 61.540 ;
        RECT 29.630 61.260 32.010 61.540 ;
        RECT 32.850 61.260 38.450 61.540 ;
        RECT 39.290 61.260 41.670 61.540 ;
        RECT 42.510 61.260 48.660 61.540 ;
        RECT 4.230 4.280 48.660 61.260 ;
        RECT 4.230 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 48.660 4.280 ;
      LAYER met3 ;
        RECT 3.990 48.640 50.820 54.565 ;
        RECT 4.400 47.240 50.820 48.640 ;
        RECT 3.990 45.240 50.820 47.240 ;
        RECT 4.400 43.840 50.820 45.240 ;
        RECT 3.990 41.840 50.820 43.840 ;
        RECT 3.990 40.440 50.420 41.840 ;
        RECT 3.990 38.440 50.820 40.440 ;
        RECT 4.400 37.040 50.420 38.440 ;
        RECT 3.990 35.040 50.820 37.040 ;
        RECT 4.400 33.640 50.420 35.040 ;
        RECT 3.990 31.640 50.820 33.640 ;
        RECT 4.400 30.240 50.420 31.640 ;
        RECT 3.990 28.240 50.820 30.240 ;
        RECT 4.400 26.840 50.420 28.240 ;
        RECT 3.990 24.840 50.820 26.840 ;
        RECT 4.400 23.440 50.420 24.840 ;
        RECT 3.990 21.440 50.820 23.440 ;
        RECT 4.400 20.040 50.420 21.440 ;
        RECT 3.990 10.715 50.820 20.040 ;
  END
END alu_8bit
END LIBRARY

