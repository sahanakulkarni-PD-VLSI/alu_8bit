VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu_8bit
  CLASS BLOCK ;
  FOREIGN alu_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 59.990 BY 70.710 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.115 10.640 15.715 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.305 10.640 27.905 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.495 10.640 40.095 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.685 10.640 52.285 57.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.155 54.520 20.755 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.710 54.520 32.310 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 42.265 54.520 43.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 53.820 54.520 55.420 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.815 10.640 12.415 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.005 10.640 24.605 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.195 10.640 36.795 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.385 10.640 48.985 57.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.855 54.520 17.455 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.410 54.520 29.010 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 38.965 54.520 40.565 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 50.520 54.520 52.120 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 55.990 23.840 59.990 24.440 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 55.990 44.240 59.990 44.840 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 66.710 39.010 70.710 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 66.710 22.910 70.710 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 55.990 27.240 59.990 27.840 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 55.990 40.840 59.990 41.440 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 66.710 35.790 70.710 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 66.710 19.690 70.710 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END b[7]
  PIN cin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END cin
  PIN cout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END cout
  PIN op[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END op[0]
  PIN op[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 55.990 34.040 59.990 34.640 ;
    END
  END op[1]
  PIN op[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 55.990 30.640 59.990 31.240 ;
    END
  END op[2]
  PIN result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END result[0]
  PIN result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 55.990 37.440 59.990 38.040 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 66.710 29.350 70.710 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END result[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 54.470 57.310 ;
      LAYER li1 ;
        RECT 5.520 10.795 54.280 57.205 ;
      LAYER met1 ;
        RECT 4.210 10.640 54.280 59.460 ;
      LAYER met2 ;
        RECT 4.230 66.430 19.130 67.050 ;
        RECT 19.970 66.430 22.350 67.050 ;
        RECT 23.190 66.430 28.790 67.050 ;
        RECT 29.630 66.430 35.230 67.050 ;
        RECT 36.070 66.430 38.450 67.050 ;
        RECT 39.290 66.430 53.730 67.050 ;
        RECT 4.230 4.280 53.730 66.430 ;
        RECT 4.230 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 53.730 4.280 ;
      LAYER met3 ;
        RECT 3.990 52.040 55.990 57.285 ;
        RECT 4.400 50.640 55.990 52.040 ;
        RECT 3.990 45.240 55.990 50.640 ;
        RECT 4.400 43.840 55.590 45.240 ;
        RECT 3.990 41.840 55.990 43.840 ;
        RECT 4.400 40.440 55.590 41.840 ;
        RECT 3.990 38.440 55.990 40.440 ;
        RECT 4.400 37.040 55.590 38.440 ;
        RECT 3.990 35.040 55.990 37.040 ;
        RECT 3.990 33.640 55.590 35.040 ;
        RECT 3.990 31.640 55.990 33.640 ;
        RECT 4.400 30.240 55.590 31.640 ;
        RECT 3.990 28.240 55.990 30.240 ;
        RECT 4.400 26.840 55.590 28.240 ;
        RECT 3.990 24.840 55.990 26.840 ;
        RECT 4.400 23.440 55.590 24.840 ;
        RECT 3.990 18.040 55.990 23.440 ;
        RECT 4.400 16.640 55.990 18.040 ;
        RECT 3.990 10.715 55.990 16.640 ;
  END
END alu_8bit
END LIBRARY

