magic
tech sky130A
magscale 1 2
timestamp 1746631653
<< nwell >>
rect 1066 2159 9882 10897
<< obsli1 >>
rect 1104 2159 9844 10897
<< obsm1 >>
rect 842 2128 9844 10928
<< metal2 >>
rect 3882 12308 3938 13108
rect 5170 12308 5226 13108
rect 5814 12308 5870 13108
rect 6458 12308 6514 13108
rect 7746 12308 7802 13108
rect 8390 12308 8446 13108
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< obsm2 >>
rect 846 12252 3826 12308
rect 3994 12252 5114 12308
rect 5282 12252 5758 12308
rect 5926 12252 6402 12308
rect 6570 12252 7690 12308
rect 7858 12252 8334 12308
rect 8502 12252 9732 12308
rect 846 856 9732 12252
rect 846 800 3182 856
rect 3350 800 3826 856
rect 3994 800 4470 856
rect 4638 800 5114 856
rect 5282 800 5758 856
rect 5926 800 7046 856
rect 7214 800 7690 856
rect 7858 800 8334 856
rect 8502 800 9732 856
<< metal3 >>
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 10164 8168 10964 8288
rect 0 7488 800 7608
rect 10164 7488 10964 7608
rect 0 6808 800 6928
rect 10164 6808 10964 6928
rect 0 6128 800 6248
rect 10164 6128 10964 6248
rect 0 5448 800 5568
rect 10164 5448 10964 5568
rect 0 4768 800 4888
rect 10164 4768 10964 4888
rect 0 4088 800 4208
rect 10164 4088 10964 4208
<< obsm3 >>
rect 798 9728 10164 10913
rect 880 9448 10164 9728
rect 798 9048 10164 9448
rect 880 8768 10164 9048
rect 798 8368 10164 8768
rect 798 8088 10084 8368
rect 798 7688 10164 8088
rect 880 7408 10084 7688
rect 798 7008 10164 7408
rect 880 6728 10084 7008
rect 798 6328 10164 6728
rect 880 6048 10084 6328
rect 798 5648 10164 6048
rect 880 5368 10084 5648
rect 798 4968 10164 5368
rect 880 4688 10084 4968
rect 798 4288 10164 4688
rect 880 4008 10084 4288
rect 798 2143 10164 4008
<< metal4 >>
rect 2036 2128 2356 10928
rect 2696 2128 3016 10928
rect 4221 2128 4541 10928
rect 4881 2128 5201 10928
rect 6406 2128 6726 10928
rect 7066 2128 7386 10928
rect 8591 2128 8911 10928
rect 9251 2128 9571 10928
<< metal5 >>
rect 1056 10288 9892 10608
rect 1056 9628 9892 9948
rect 1056 8113 9892 8433
rect 1056 7453 9892 7773
rect 1056 5938 9892 6258
rect 1056 5278 9892 5598
rect 1056 3763 9892 4083
rect 1056 3103 9892 3423
<< labels >>
rlabel metal4 s 2696 2128 3016 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4881 2128 5201 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7066 2128 7386 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9251 2128 9571 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3763 9892 4083 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5938 9892 6258 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8113 9892 8433 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 10288 9892 10608 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2036 2128 2356 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4221 2128 4541 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6406 2128 6726 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8591 2128 8911 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3103 9892 3423 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5278 9892 5598 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7453 9892 7773 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 9628 9892 9948 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 8390 0 8446 800 6 a[0]
port 3 nsew signal input
rlabel metal3 s 10164 4768 10964 4888 6 a[1]
port 4 nsew signal input
rlabel metal2 s 7746 12308 7802 13108 6 a[2]
port 5 nsew signal input
rlabel metal2 s 6458 12308 6514 13108 6 a[3]
port 6 nsew signal input
rlabel metal2 s 3882 12308 3938 13108 6 a[4]
port 7 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 a[5]
port 8 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 a[6]
port 9 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 a[7]
port 10 nsew signal input
rlabel metal3 s 10164 4088 10964 4208 6 b[0]
port 11 nsew signal input
rlabel metal3 s 10164 5448 10964 5568 6 b[1]
port 12 nsew signal input
rlabel metal2 s 8390 12308 8446 13108 6 b[2]
port 13 nsew signal input
rlabel metal2 s 5814 12308 5870 13108 6 b[3]
port 14 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 b[4]
port 15 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 b[5]
port 16 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 b[6]
port 17 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 b[7]
port 18 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 cin
port 19 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 cout
port 20 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 op[0]
port 21 nsew signal input
rlabel metal3 s 10164 6808 10964 6928 6 op[1]
port 22 nsew signal input
rlabel metal3 s 10164 8168 10964 8288 6 op[2]
port 23 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 result[0]
port 24 nsew signal output
rlabel metal3 s 10164 6128 10964 6248 6 result[1]
port 25 nsew signal output
rlabel metal3 s 10164 7488 10964 7608 6 result[2]
port 26 nsew signal output
rlabel metal2 s 5170 12308 5226 13108 6 result[3]
port 27 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 result[4]
port 28 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 result[5]
port 29 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 result[6]
port 30 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 result[7]
port 31 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 10964 13108
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 731162
string GDS_FILE /openlane/designs/alu_8bit/runs/RUN_2025.05.07_15.24.49/results/signoff/alu_8bit.magic.gds
string GDS_START 321248
<< end >>

