magic
tech sky130A
magscale 1 2
timestamp 1746639707
<< checkpaint >>
rect -3932 -3932 14133 16277
<< viali >>
rect 3525 9605 3559 9639
rect 4353 9605 4387 9639
rect 1409 9537 1443 9571
rect 1961 9537 1995 9571
rect 2053 9537 2087 9571
rect 3065 9537 3099 9571
rect 4077 9537 4111 9571
rect 4721 9537 4755 9571
rect 5089 9537 5123 9571
rect 5457 9537 5491 9571
rect 6469 9537 6503 9571
rect 6745 9537 6779 9571
rect 7205 9537 7239 9571
rect 7481 9537 7515 9571
rect 7665 9537 7699 9571
rect 7757 9537 7791 9571
rect 8033 9537 8067 9571
rect 8217 9537 8251 9571
rect 8677 9537 8711 9571
rect 5273 9469 5307 9503
rect 5549 9469 5583 9503
rect 6377 9469 6411 9503
rect 6929 9469 6963 9503
rect 4261 9401 4295 9435
rect 5089 9401 5123 9435
rect 7849 9401 7883 9435
rect 8493 9401 8527 9435
rect 1593 9333 1627 9367
rect 1777 9333 1811 9367
rect 2237 9333 2271 9367
rect 3157 9333 3191 9367
rect 3433 9333 3467 9367
rect 6009 9333 6043 9367
rect 7021 9333 7055 9367
rect 7573 9333 7607 9367
rect 8033 9333 8067 9367
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 2973 9061 3007 9095
rect 1593 8993 1627 9027
rect 2237 8993 2271 9027
rect 3617 8993 3651 9027
rect 4997 8993 5031 9027
rect 6653 8993 6687 9027
rect 7113 8993 7147 9027
rect 8585 8993 8619 9027
rect 1777 8925 1811 8959
rect 1869 8925 1903 8959
rect 2329 8925 2363 8959
rect 3801 8925 3835 8959
rect 4261 8925 4295 8959
rect 4629 8925 4663 8959
rect 4813 8925 4847 8959
rect 5365 8925 5399 8959
rect 5549 8925 5583 8959
rect 6285 8925 6319 8959
rect 7297 8925 7331 8959
rect 7665 8925 7699 8959
rect 7849 8925 7883 8959
rect 8125 8925 8159 8959
rect 8427 8925 8461 8959
rect 2605 8857 2639 8891
rect 2821 8857 2855 8891
rect 3985 8857 4019 8891
rect 6101 8857 6135 8891
rect 7941 8857 7975 8891
rect 8217 8857 8251 8891
rect 8309 8857 8343 8891
rect 1593 8789 1627 8823
rect 1961 8789 1995 8823
rect 3157 8789 3191 8823
rect 4169 8789 4203 8823
rect 4629 8789 4663 8823
rect 6469 8789 6503 8823
rect 2897 8585 2931 8619
rect 4813 8585 4847 8619
rect 5181 8585 5215 8619
rect 8033 8585 8067 8619
rect 2237 8517 2271 8551
rect 2697 8517 2731 8551
rect 3249 8517 3283 8551
rect 5641 8517 5675 8551
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2145 8449 2179 8483
rect 2421 8449 2455 8483
rect 2513 8449 2547 8483
rect 3157 8449 3191 8483
rect 3433 8449 3467 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 4077 8449 4111 8483
rect 4169 8449 4203 8483
rect 4629 8449 4663 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 5457 8449 5491 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 6653 8449 6687 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 8493 8449 8527 8483
rect 3617 8381 3651 8415
rect 6377 8381 6411 8415
rect 8217 8381 8251 8415
rect 8309 8381 8343 8415
rect 8401 8381 8435 8415
rect 1501 8313 1535 8347
rect 2053 8313 2087 8347
rect 5273 8313 5307 8347
rect 6101 8313 6135 8347
rect 2237 8245 2271 8279
rect 2881 8245 2915 8279
rect 3065 8245 3099 8279
rect 4353 8245 4387 8279
rect 5825 8245 5859 8279
rect 7481 8245 7515 8279
rect 4629 8041 4663 8075
rect 7205 8041 7239 8075
rect 3985 7905 4019 7939
rect 4077 7905 4111 7939
rect 6009 7905 6043 7939
rect 7481 7905 7515 7939
rect 7758 7905 7792 7939
rect 2237 7837 2271 7871
rect 2329 7837 2363 7871
rect 2789 7837 2823 7871
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 4905 7837 4939 7871
rect 5273 7837 5307 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 7665 7837 7699 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 8401 7837 8435 7871
rect 1777 7769 1811 7803
rect 1961 7769 1995 7803
rect 2605 7769 2639 7803
rect 2697 7769 2731 7803
rect 4997 7769 5031 7803
rect 5135 7769 5169 7803
rect 5917 7769 5951 7803
rect 1593 7701 1627 7735
rect 2053 7701 2087 7735
rect 2973 7701 3007 7735
rect 4353 7701 4387 7735
rect 5365 7701 5399 7735
rect 7297 7701 7331 7735
rect 8125 7701 8159 7735
rect 8585 7701 8619 7735
rect 2237 7497 2271 7531
rect 4905 7497 4939 7531
rect 7757 7497 7791 7531
rect 1731 7429 1765 7463
rect 1961 7429 1995 7463
rect 4537 7429 4571 7463
rect 6561 7429 6595 7463
rect 8033 7429 8067 7463
rect 1593 7361 1627 7395
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 4721 7361 4755 7395
rect 5457 7361 5491 7395
rect 6009 7361 6043 7395
rect 6653 7361 6687 7395
rect 6745 7361 6779 7395
rect 6837 7361 6871 7395
rect 7021 7361 7055 7395
rect 7113 7361 7147 7395
rect 7292 7361 7326 7395
rect 7389 7361 7423 7395
rect 7481 7361 7515 7395
rect 8585 7361 8619 7395
rect 5273 7293 5307 7327
rect 7021 7157 7055 7191
rect 3433 6953 3467 6987
rect 4537 6953 4571 6987
rect 7297 6953 7331 6987
rect 5733 6885 5767 6919
rect 7757 6885 7791 6919
rect 5365 6817 5399 6851
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 5181 6749 5215 6783
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 6926 6749 6960 6783
rect 7389 6749 7423 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 8493 6749 8527 6783
rect 2329 6681 2363 6715
rect 2513 6681 2547 6715
rect 3249 6681 3283 6715
rect 4505 6681 4539 6715
rect 4721 6681 4755 6715
rect 4997 6681 5031 6715
rect 5457 6681 5491 6715
rect 8677 6681 8711 6715
rect 1501 6613 1535 6647
rect 1777 6613 1811 6647
rect 2145 6613 2179 6647
rect 3454 6613 3488 6647
rect 3617 6613 3651 6647
rect 3801 6613 3835 6647
rect 4353 6613 4387 6647
rect 5917 6613 5951 6647
rect 6377 6613 6411 6647
rect 6745 6613 6779 6647
rect 6929 6613 6963 6647
rect 2973 6409 3007 6443
rect 6101 6409 6135 6443
rect 1777 6341 1811 6375
rect 1961 6341 1995 6375
rect 3065 6341 3099 6375
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2789 6273 2823 6307
rect 2973 6273 3007 6307
rect 3249 6273 3283 6307
rect 4077 6273 4111 6307
rect 4445 6273 4479 6307
rect 4905 6273 4939 6307
rect 5273 6273 5307 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 5825 6273 5859 6307
rect 5917 6273 5951 6307
rect 6469 6273 6503 6307
rect 6561 6273 6595 6307
rect 7297 6273 7331 6307
rect 8585 6273 8619 6307
rect 2605 6205 2639 6239
rect 2697 6205 2731 6239
rect 3433 6205 3467 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 3985 6205 4019 6239
rect 6653 6205 6687 6239
rect 8033 6205 8067 6239
rect 5457 6137 5491 6171
rect 1593 6069 1627 6103
rect 2053 6069 2087 6103
rect 5089 6069 5123 6103
rect 7113 6069 7147 6103
rect 7757 6069 7791 6103
rect 1593 5865 1627 5899
rect 3893 5865 3927 5899
rect 8493 5865 8527 5899
rect 1685 5729 1719 5763
rect 2513 5729 2547 5763
rect 4261 5729 4295 5763
rect 4353 5729 4387 5763
rect 5273 5729 5307 5763
rect 7021 5729 7055 5763
rect 8125 5729 8159 5763
rect 8217 5729 8251 5763
rect 8401 5729 8435 5763
rect 1409 5661 1443 5695
rect 2053 5661 2087 5695
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 3249 5661 3283 5695
rect 3801 5661 3835 5695
rect 4445 5661 4479 5695
rect 4629 5661 4663 5695
rect 4813 5661 4847 5695
rect 5641 5661 5675 5695
rect 6561 5661 6595 5695
rect 6653 5661 6687 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8033 5661 8067 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 1823 5593 1857 5627
rect 1961 5593 1995 5627
rect 4997 5593 5031 5627
rect 5457 5593 5491 5627
rect 5917 5593 5951 5627
rect 6101 5593 6135 5627
rect 6929 5593 6963 5627
rect 3341 5525 3375 5559
rect 5089 5525 5123 5559
rect 5733 5525 5767 5559
rect 6377 5525 6411 5559
rect 7205 5525 7239 5559
rect 1961 5321 1995 5355
rect 4261 5321 4295 5355
rect 6377 5321 6411 5355
rect 4813 5253 4847 5287
rect 5963 5253 5997 5287
rect 1685 5185 1719 5219
rect 1777 5185 1811 5219
rect 2237 5185 2271 5219
rect 3341 5185 3375 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 3709 5185 3743 5219
rect 4169 5185 4203 5219
rect 4537 5185 4571 5219
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 5733 5185 5767 5219
rect 5825 5185 5859 5219
rect 6101 5185 6135 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 7297 5185 7331 5219
rect 7665 5185 7699 5219
rect 4445 5117 4479 5151
rect 4905 5117 4939 5151
rect 2053 5049 2087 5083
rect 7389 5049 7423 5083
rect 1501 4981 1535 5015
rect 3157 4981 3191 5015
rect 3985 4981 4019 5015
rect 5365 4981 5399 5015
rect 6745 4777 6779 4811
rect 8493 4777 8527 4811
rect 5273 4709 5307 4743
rect 7481 4709 7515 4743
rect 2237 4641 2271 4675
rect 2605 4641 2639 4675
rect 4261 4641 4295 4675
rect 5733 4641 5767 4675
rect 6285 4641 6319 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 1777 4573 1811 4607
rect 2329 4573 2363 4607
rect 2697 4573 2731 4607
rect 3801 4573 3835 4607
rect 4353 4573 4387 4607
rect 6009 4573 6043 4607
rect 7941 4573 7975 4607
rect 1961 4505 1995 4539
rect 5825 4505 5859 4539
rect 1593 4437 1627 4471
rect 2053 4437 2087 4471
rect 3985 4437 4019 4471
rect 2237 4233 2271 4267
rect 2897 4233 2931 4267
rect 4261 4233 4295 4267
rect 4813 4233 4847 4267
rect 6377 4233 6411 4267
rect 7021 4233 7055 4267
rect 7573 4233 7607 4267
rect 1751 4165 1785 4199
rect 2697 4165 2731 4199
rect 6745 4165 6779 4199
rect 1593 4097 1627 4131
rect 1869 4097 1903 4131
rect 1961 4097 1995 4131
rect 2053 4097 2087 4131
rect 4077 4097 4111 4131
rect 4721 4097 4755 4131
rect 5089 4097 5123 4131
rect 5273 4097 5307 4131
rect 5641 4097 5675 4131
rect 5733 4097 5767 4131
rect 5917 4097 5951 4131
rect 6193 4097 6227 4131
rect 6561 4097 6595 4131
rect 6837 4097 6871 4131
rect 7021 4097 7055 4131
rect 7297 4097 7331 4131
rect 7757 4097 7791 4131
rect 7941 4097 7975 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 3801 4029 3835 4063
rect 4997 4029 5031 4063
rect 5181 4029 5215 4063
rect 7113 4029 7147 4063
rect 7665 4029 7699 4063
rect 3065 3961 3099 3995
rect 3893 3961 3927 3995
rect 6009 3961 6043 3995
rect 8585 3961 8619 3995
rect 2881 3893 2915 3927
rect 3985 3893 4019 3927
rect 5457 3893 5491 3927
rect 5825 3893 5859 3927
rect 1869 3689 1903 3723
rect 2145 3689 2179 3723
rect 2789 3689 2823 3723
rect 4169 3689 4203 3723
rect 5273 3689 5307 3723
rect 1593 3621 1627 3655
rect 3157 3621 3191 3655
rect 4353 3621 4387 3655
rect 6561 3621 6595 3655
rect 1961 3553 1995 3587
rect 4813 3553 4847 3587
rect 5181 3553 5215 3587
rect 5917 3553 5951 3587
rect 8401 3553 8435 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 1777 3485 1811 3519
rect 2053 3485 2087 3519
rect 2237 3485 2271 3519
rect 2421 3485 2455 3519
rect 2881 3485 2915 3519
rect 3341 3485 3375 3519
rect 3617 3485 3651 3519
rect 4629 3485 4663 3519
rect 4905 3485 4939 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6193 3485 6227 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7297 3485 7331 3519
rect 7573 3485 7607 3519
rect 7849 3485 7883 3519
rect 8042 3485 8076 3519
rect 2605 3417 2639 3451
rect 3985 3417 4019 3451
rect 4185 3417 4219 3451
rect 4445 3417 4479 3451
rect 6101 3417 6135 3451
rect 2973 3349 3007 3383
rect 3433 3349 3467 3383
rect 5457 3349 5491 3383
rect 5641 3349 5675 3383
rect 6837 3349 6871 3383
rect 1961 3145 1995 3179
rect 3525 3145 3559 3179
rect 4169 3145 4203 3179
rect 5089 3145 5123 3179
rect 8125 3145 8159 3179
rect 8401 3145 8435 3179
rect 2053 3077 2087 3111
rect 2269 3077 2303 3111
rect 3801 3077 3835 3111
rect 4017 3077 4051 3111
rect 4997 3077 5031 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 2605 3009 2639 3043
rect 2789 3009 2823 3043
rect 2881 3009 2915 3043
rect 3157 3009 3191 3043
rect 3341 3009 3375 3043
rect 3617 3009 3651 3043
rect 4261 3009 4295 3043
rect 4537 3009 4571 3043
rect 5457 3009 5491 3043
rect 5549 3009 5583 3043
rect 6193 3009 6227 3043
rect 6653 3009 6687 3043
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 7757 3009 7791 3043
rect 8125 3009 8159 3043
rect 8309 3009 8343 3043
rect 8585 3009 8619 3043
rect 1685 2941 1719 2975
rect 6469 2941 6503 2975
rect 7021 2941 7055 2975
rect 7481 2941 7515 2975
rect 7573 2941 7607 2975
rect 2421 2873 2455 2907
rect 4353 2873 4387 2907
rect 6929 2873 6963 2907
rect 1685 2805 1719 2839
rect 2237 2805 2271 2839
rect 3065 2805 3099 2839
rect 3985 2805 4019 2839
rect 5733 2805 5767 2839
rect 6009 2805 6043 2839
rect 7113 2805 7147 2839
rect 1961 2601 1995 2635
rect 3341 2601 3375 2635
rect 6377 2601 6411 2635
rect 7205 2601 7239 2635
rect 7665 2601 7699 2635
rect 8493 2601 8527 2635
rect 2605 2533 2639 2567
rect 3157 2533 3191 2567
rect 6745 2533 6779 2567
rect 7757 2533 7791 2567
rect 6837 2465 6871 2499
rect 8677 2465 8711 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 2237 2397 2271 2431
rect 2513 2397 2547 2431
rect 2697 2397 2731 2431
rect 2789 2397 2823 2431
rect 3065 2397 3099 2431
rect 3249 2397 3283 2431
rect 3341 2397 3375 2431
rect 3525 2397 3559 2431
rect 3617 2397 3651 2431
rect 4077 2397 4111 2431
rect 5457 2397 5491 2431
rect 5825 2397 5859 2431
rect 6561 2397 6595 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7389 2397 7423 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 1961 2329 1995 2363
rect 4445 2329 4479 2363
rect 5089 2329 5123 2363
rect 6009 2329 6043 2363
rect 6193 2329 6227 2363
rect 8125 2329 8159 2363
rect 1593 2261 1627 2295
rect 1869 2261 1903 2295
rect 2145 2261 2179 2295
rect 2973 2261 3007 2295
<< metal1 >>
rect 1104 9818 9016 9840
rect 1104 9766 2599 9818
rect 2651 9766 2663 9818
rect 2715 9766 2727 9818
rect 2779 9766 2791 9818
rect 2843 9766 2855 9818
rect 2907 9766 4577 9818
rect 4629 9766 4641 9818
rect 4693 9766 4705 9818
rect 4757 9766 4769 9818
rect 4821 9766 4833 9818
rect 4885 9766 6555 9818
rect 6607 9766 6619 9818
rect 6671 9766 6683 9818
rect 6735 9766 6747 9818
rect 6799 9766 6811 9818
rect 6863 9766 8533 9818
rect 8585 9766 8597 9818
rect 8649 9766 8661 9818
rect 8713 9766 8725 9818
rect 8777 9766 8789 9818
rect 8841 9766 9016 9818
rect 1104 9744 9016 9766
rect 1026 9596 1032 9648
rect 1084 9636 1090 9648
rect 1084 9608 2084 9636
rect 1084 9596 1090 9608
rect 1394 9528 1400 9580
rect 1452 9528 1458 9580
rect 2056 9577 2084 9608
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3513 9639 3571 9645
rect 3513 9636 3525 9639
rect 3016 9608 3525 9636
rect 3016 9596 3022 9608
rect 3513 9605 3525 9608
rect 3559 9605 3571 9639
rect 3513 9599 3571 9605
rect 4341 9639 4399 9645
rect 4341 9605 4353 9639
rect 4387 9636 4399 9639
rect 4430 9636 4436 9648
rect 4387 9608 4436 9636
rect 4387 9605 4399 9608
rect 4341 9599 4399 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 5166 9636 5172 9648
rect 4632 9608 5172 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 1964 9500 1992 9531
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3786 9568 3792 9580
rect 3108 9540 3792 9568
rect 3108 9528 3114 9540
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4632 9568 4660 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 5868 9608 7236 9636
rect 5868 9596 5874 9608
rect 4111 9540 4660 9568
rect 4709 9571 4767 9577
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4982 9568 4988 9580
rect 4755 9540 4988 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5074 9528 5080 9580
rect 5132 9528 5138 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 6457 9571 6515 9577
rect 6457 9568 6469 9571
rect 5491 9540 6469 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 6457 9537 6469 9540
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7208 9577 7236 9608
rect 7484 9608 7788 9636
rect 7484 9577 7512 9608
rect 7760 9580 7788 9608
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 7616 9540 7665 9568
rect 7616 9528 7622 9540
rect 7653 9537 7665 9540
rect 7699 9537 7711 9571
rect 7653 9531 7711 9537
rect 2406 9500 2412 9512
rect 1964 9472 2412 9500
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 5092 9500 5120 9528
rect 4264 9472 5120 9500
rect 4264 9441 4292 9472
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5316 9472 5549 9500
rect 5316 9460 5322 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6696 9472 6929 9500
rect 6696 9460 6702 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 7668 9500 7696 9531
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7800 9540 8033 9568
rect 7800 9528 7806 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 8938 9568 8944 9580
rect 8711 9540 8944 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 8220 9500 8248 9531
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 7668 9472 8524 9500
rect 6917 9463 6975 9469
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9401 4307 9435
rect 4249 9395 4307 9401
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4396 9404 5089 9432
rect 4396 9392 4402 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 5077 9395 5135 9401
rect 7837 9435 7895 9441
rect 7837 9401 7849 9435
rect 7883 9432 7895 9435
rect 8386 9432 8392 9444
rect 7883 9404 8392 9432
rect 7883 9401 7895 9404
rect 7837 9395 7895 9401
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8496 9441 8524 9472
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9401 8539 9435
rect 8481 9395 8539 9401
rect 1578 9324 1584 9376
rect 1636 9324 1642 9376
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 1765 9367 1823 9373
rect 1765 9364 1777 9367
rect 1728 9336 1777 9364
rect 1728 9324 1734 9336
rect 1765 9333 1777 9336
rect 1811 9333 1823 9367
rect 1765 9327 1823 9333
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2590 9364 2596 9376
rect 2271 9336 2596 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 3142 9324 3148 9376
rect 3200 9324 3206 9376
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 3602 9364 3608 9376
rect 3467 9336 3608 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5684 9336 6009 9364
rect 5684 9324 5690 9336
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 5997 9327 6055 9333
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6788 9336 7021 9364
rect 6788 9324 6794 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7432 9336 7573 9364
rect 7432 9324 7438 9336
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 7561 9327 7619 9333
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 8294 9364 8300 9376
rect 8067 9336 8300 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 1104 9274 9016 9296
rect 1104 9222 1939 9274
rect 1991 9222 2003 9274
rect 2055 9222 2067 9274
rect 2119 9222 2131 9274
rect 2183 9222 2195 9274
rect 2247 9222 3917 9274
rect 3969 9222 3981 9274
rect 4033 9222 4045 9274
rect 4097 9222 4109 9274
rect 4161 9222 4173 9274
rect 4225 9222 5895 9274
rect 5947 9222 5959 9274
rect 6011 9222 6023 9274
rect 6075 9222 6087 9274
rect 6139 9222 6151 9274
rect 6203 9222 7873 9274
rect 7925 9222 7937 9274
rect 7989 9222 8001 9274
rect 8053 9222 8065 9274
rect 8117 9222 8129 9274
rect 8181 9222 9016 9274
rect 1104 9200 9016 9222
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9129 2375 9163
rect 2317 9123 2375 9129
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3234 9160 3240 9172
rect 2823 9132 3240 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 1854 9052 1860 9104
rect 1912 9092 1918 9104
rect 2332 9092 2360 9123
rect 3234 9120 3240 9132
rect 3292 9160 3298 9172
rect 4338 9160 4344 9172
rect 3292 9132 4344 9160
rect 3292 9120 3298 9132
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 4540 9132 5304 9160
rect 2961 9095 3019 9101
rect 2961 9092 2973 9095
rect 1912 9064 2973 9092
rect 1912 9052 1918 9064
rect 2961 9061 2973 9064
rect 3007 9092 3019 9095
rect 3510 9092 3516 9104
rect 3007 9064 3516 9092
rect 3007 9061 3019 9064
rect 2961 9055 3019 9061
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 4540 9092 4568 9132
rect 5166 9092 5172 9104
rect 4172 9064 4568 9092
rect 4632 9064 5172 9092
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 1946 9024 1952 9036
rect 1636 8996 1952 9024
rect 1636 8984 1642 8996
rect 1946 8984 1952 8996
rect 2004 9024 2010 9036
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 2004 8996 2237 9024
rect 2004 8984 2010 8996
rect 2225 8993 2237 8996
rect 2271 9024 2283 9027
rect 3050 9024 3056 9036
rect 2271 8996 3056 9024
rect 2271 8993 2283 8996
rect 2225 8987 2283 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 3602 8984 3608 9036
rect 3660 8984 3666 9036
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 1780 8888 1808 8919
rect 1854 8916 1860 8968
rect 1912 8916 1918 8968
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 3418 8956 3424 8968
rect 2317 8919 2375 8925
rect 2746 8928 3424 8956
rect 2222 8888 2228 8900
rect 1780 8860 2228 8888
rect 2222 8848 2228 8860
rect 2280 8888 2286 8900
rect 2332 8888 2360 8919
rect 2280 8860 2360 8888
rect 2280 8848 2286 8860
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 2746 8888 2774 8928
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 2648 8860 2774 8888
rect 2809 8891 2867 8897
rect 2648 8848 2654 8860
rect 2809 8857 2821 8891
rect 2855 8888 2867 8891
rect 3326 8888 3332 8900
rect 2855 8860 3332 8888
rect 2855 8857 2867 8860
rect 2809 8851 2867 8857
rect 3326 8848 3332 8860
rect 3384 8888 3390 8900
rect 3620 8888 3648 8984
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 4172 8956 4200 9064
rect 3896 8928 4200 8956
rect 4249 8959 4307 8965
rect 3384 8860 3648 8888
rect 3384 8848 3390 8860
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 3896 8888 3924 8928
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4430 8956 4436 8968
rect 4295 8928 4436 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4632 8965 4660 9064
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5276 9092 5304 9132
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 7616 9132 8248 9160
rect 7616 9120 7622 9132
rect 6362 9092 6368 9104
rect 5276 9064 6368 9092
rect 6362 9052 6368 9064
rect 6420 9092 6426 9104
rect 6420 9064 7144 9092
rect 6420 9052 6426 9064
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5258 9024 5264 9036
rect 5031 8996 5264 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 6638 9024 6644 9036
rect 5368 8996 6644 9024
rect 5368 8965 5396 8996
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 7116 9033 7144 9064
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8220 9024 8248 9132
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 8076 8996 8156 9024
rect 8220 8996 8585 9024
rect 8076 8984 8082 8996
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8956 4859 8959
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 4847 8928 5365 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 6273 8959 6331 8965
rect 6273 8956 6285 8959
rect 5592 8928 6285 8956
rect 5592 8916 5598 8928
rect 6273 8925 6285 8928
rect 6319 8956 6331 8959
rect 6730 8956 6736 8968
rect 6319 8928 6736 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 3752 8860 3924 8888
rect 3973 8891 4031 8897
rect 3752 8848 3758 8860
rect 3973 8857 3985 8891
rect 4019 8857 4031 8891
rect 3973 8851 4031 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1762 8820 1768 8832
rect 1627 8792 1768 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 1854 8780 1860 8832
rect 1912 8820 1918 8832
rect 1949 8823 2007 8829
rect 1949 8820 1961 8823
rect 1912 8792 1961 8820
rect 1912 8780 1918 8792
rect 1949 8789 1961 8792
rect 1995 8789 2007 8823
rect 1949 8783 2007 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 3108 8792 3157 8820
rect 3108 8780 3114 8792
rect 3145 8789 3157 8792
rect 3191 8789 3203 8823
rect 3145 8783 3203 8789
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 3988 8820 4016 8851
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 6089 8891 6147 8897
rect 6089 8888 6101 8891
rect 5132 8860 6101 8888
rect 5132 8848 5138 8860
rect 6089 8857 6101 8860
rect 6135 8857 6147 8891
rect 7300 8888 7328 8919
rect 7650 8916 7656 8968
rect 7708 8916 7714 8968
rect 8128 8965 8156 8996
rect 8573 8993 8585 8996
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8113 8959 8171 8965
rect 7883 8928 8064 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 7929 8891 7987 8897
rect 7929 8888 7941 8891
rect 7300 8860 7941 8888
rect 6089 8851 6147 8857
rect 7929 8857 7941 8860
rect 7975 8857 7987 8891
rect 7929 8851 7987 8857
rect 3476 8792 4016 8820
rect 4157 8823 4215 8829
rect 3476 8780 3482 8792
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4246 8820 4252 8832
rect 4203 8792 4252 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4617 8823 4675 8829
rect 4617 8789 4629 8823
rect 4663 8820 4675 8823
rect 5994 8820 6000 8832
rect 4663 8792 6000 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 6236 8792 6469 8820
rect 6236 8780 6242 8792
rect 6457 8789 6469 8792
rect 6503 8789 6515 8823
rect 8036 8820 8064 8928
rect 8113 8925 8125 8959
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8386 8916 8392 8968
rect 8444 8965 8450 8968
rect 8444 8959 8473 8965
rect 8461 8925 8473 8959
rect 8444 8919 8473 8925
rect 8444 8916 8450 8919
rect 8202 8848 8208 8900
rect 8260 8848 8266 8900
rect 8297 8891 8355 8897
rect 8297 8857 8309 8891
rect 8343 8888 8355 8891
rect 9030 8888 9036 8900
rect 8343 8860 9036 8888
rect 8343 8857 8355 8860
rect 8297 8851 8355 8857
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 8386 8820 8392 8832
rect 8036 8792 8392 8820
rect 6457 8783 6515 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 1104 8730 9016 8752
rect 1104 8678 2599 8730
rect 2651 8678 2663 8730
rect 2715 8678 2727 8730
rect 2779 8678 2791 8730
rect 2843 8678 2855 8730
rect 2907 8678 4577 8730
rect 4629 8678 4641 8730
rect 4693 8678 4705 8730
rect 4757 8678 4769 8730
rect 4821 8678 4833 8730
rect 4885 8678 6555 8730
rect 6607 8678 6619 8730
rect 6671 8678 6683 8730
rect 6735 8678 6747 8730
rect 6799 8678 6811 8730
rect 6863 8678 8533 8730
rect 8585 8678 8597 8730
rect 8649 8678 8661 8730
rect 8713 8678 8725 8730
rect 8777 8678 8789 8730
rect 8841 8678 9016 8730
rect 1104 8656 9016 8678
rect 2498 8576 2504 8628
rect 2556 8576 2562 8628
rect 2866 8576 2872 8628
rect 2924 8625 2930 8628
rect 2924 8619 2943 8625
rect 2931 8585 2943 8619
rect 2924 8579 2943 8585
rect 2924 8576 2930 8579
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4801 8619 4859 8625
rect 3200 8588 4108 8616
rect 3200 8576 3206 8588
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8548 2283 8551
rect 2516 8548 2544 8576
rect 2271 8520 2544 8548
rect 2271 8517 2283 8520
rect 2225 8511 2283 8517
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1946 8440 1952 8492
rect 2004 8440 2010 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2240 8480 2268 8511
rect 2682 8508 2688 8560
rect 2740 8508 2746 8560
rect 3234 8508 3240 8560
rect 3292 8508 3298 8560
rect 3694 8508 3700 8560
rect 3752 8548 3758 8560
rect 4080 8548 4108 8588
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 4982 8616 4988 8628
rect 4847 8588 4988 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 5442 8616 5448 8628
rect 5224 8588 5448 8616
rect 5224 8576 5230 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7708 8588 8033 8616
rect 7708 8576 7714 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 5534 8548 5540 8560
rect 3752 8520 3924 8548
rect 4080 8520 4200 8548
rect 3752 8508 3758 8520
rect 2179 8452 2268 8480
rect 2409 8483 2467 8489
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 3050 8480 3056 8492
rect 2547 8452 3056 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2424 8412 2452 8443
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3142 8440 3148 8492
rect 3200 8440 3206 8492
rect 2682 8412 2688 8424
rect 2424 8384 2688 8412
rect 2682 8372 2688 8384
rect 2740 8412 2746 8424
rect 3252 8412 3280 8508
rect 3418 8440 3424 8492
rect 3476 8440 3482 8492
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3896 8489 3924 8520
rect 4172 8489 4200 8520
rect 5184 8520 5540 8548
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 3568 8452 3801 8480
rect 3568 8440 3574 8452
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 2740 8384 3280 8412
rect 3605 8415 3663 8421
rect 2740 8372 2746 8384
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 4080 8412 4108 8443
rect 4614 8440 4620 8492
rect 4672 8440 4678 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5074 8480 5080 8492
rect 5031 8452 5080 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5184 8489 5212 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 5626 8508 5632 8560
rect 5684 8548 5690 8560
rect 5684 8520 5856 8548
rect 5684 8508 5690 8520
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5491 8452 5733 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 3651 8384 4108 8412
rect 5092 8412 5120 8440
rect 5460 8412 5488 8443
rect 5092 8384 5488 8412
rect 5828 8412 5856 8520
rect 5920 8520 6684 8548
rect 5920 8489 5948 8520
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6656 8489 6684 8520
rect 8294 8508 8300 8560
rect 8352 8508 8358 8560
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7800 8452 7849 8480
rect 7800 8440 7806 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 8312 8480 8340 8508
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8312 8452 8493 8480
rect 7837 8443 7895 8449
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5828 8384 6377 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 8076 8384 8217 8412
rect 8076 8372 8082 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 2314 8344 2320 8356
rect 2087 8316 2320 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 2314 8304 2320 8316
rect 2372 8344 2378 8356
rect 2372 8316 2774 8344
rect 2372 8304 2378 8316
rect 2222 8236 2228 8288
rect 2280 8236 2286 8288
rect 2746 8276 2774 8316
rect 2958 8304 2964 8356
rect 3016 8344 3022 8356
rect 3016 8316 4476 8344
rect 3016 8304 3022 8316
rect 2869 8279 2927 8285
rect 2869 8276 2881 8279
rect 2746 8248 2881 8276
rect 2869 8245 2881 8248
rect 2915 8245 2927 8279
rect 2869 8239 2927 8245
rect 3050 8236 3056 8288
rect 3108 8236 3114 8288
rect 4338 8236 4344 8288
rect 4396 8236 4402 8288
rect 4448 8276 4476 8316
rect 4890 8304 4896 8356
rect 4948 8344 4954 8356
rect 5261 8347 5319 8353
rect 5261 8344 5273 8347
rect 4948 8316 5273 8344
rect 4948 8304 4954 8316
rect 5261 8313 5273 8316
rect 5307 8313 5319 8347
rect 6089 8347 6147 8353
rect 6089 8344 6101 8347
rect 5261 8307 5319 8313
rect 5368 8316 6101 8344
rect 5368 8276 5396 8316
rect 6089 8313 6101 8316
rect 6135 8313 6147 8347
rect 8220 8344 8248 8375
rect 8294 8372 8300 8424
rect 8352 8372 8358 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8412 8447 8415
rect 9030 8412 9036 8424
rect 8435 8384 9036 8412
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 9122 8344 9128 8356
rect 8220 8316 9128 8344
rect 6089 8307 6147 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 4448 8248 5396 8276
rect 5810 8236 5816 8288
rect 5868 8236 5874 8288
rect 7466 8236 7472 8288
rect 7524 8236 7530 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8110 8276 8116 8288
rect 7708 8248 8116 8276
rect 7708 8236 7714 8248
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 1104 8186 9016 8208
rect 1104 8134 1939 8186
rect 1991 8134 2003 8186
rect 2055 8134 2067 8186
rect 2119 8134 2131 8186
rect 2183 8134 2195 8186
rect 2247 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 5895 8186
rect 5947 8134 5959 8186
rect 6011 8134 6023 8186
rect 6075 8134 6087 8186
rect 6139 8134 6151 8186
rect 6203 8134 7873 8186
rect 7925 8134 7937 8186
rect 7989 8134 8001 8186
rect 8053 8134 8065 8186
rect 8117 8134 8129 8186
rect 8181 8134 9016 8186
rect 1104 8112 9016 8134
rect 4614 8032 4620 8084
rect 4672 8032 4678 8084
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7742 8072 7748 8084
rect 7239 8044 7748 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 7484 7976 7972 8004
rect 7484 7948 7512 7976
rect 1302 7896 1308 7948
rect 1360 7936 1366 7948
rect 1360 7908 2820 7936
rect 1360 7896 1366 7908
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 2792 7877 2820 7908
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 3973 7939 4031 7945
rect 3973 7936 3985 7939
rect 3108 7908 3985 7936
rect 3108 7896 3114 7908
rect 3973 7905 3985 7908
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4430 7936 4436 7948
rect 4111 7908 4436 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 5810 7936 5816 7948
rect 4816 7908 5816 7936
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 4246 7828 4252 7880
rect 4304 7828 4310 7880
rect 4816 7877 4844 7908
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7936 6055 7939
rect 6270 7936 6276 7948
rect 6043 7908 6276 7936
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7374 7936 7380 7948
rect 6972 7908 7380 7936
rect 6972 7896 6978 7908
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 7466 7896 7472 7948
rect 7524 7896 7530 7948
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 1394 7760 1400 7812
rect 1452 7800 1458 7812
rect 1765 7803 1823 7809
rect 1765 7800 1777 7803
rect 1452 7772 1777 7800
rect 1452 7760 1458 7772
rect 1765 7769 1777 7772
rect 1811 7769 1823 7803
rect 1765 7763 1823 7769
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7800 2007 7803
rect 2332 7800 2360 7828
rect 1995 7772 2360 7800
rect 1995 7769 2007 7772
rect 1949 7763 2007 7769
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 2593 7803 2651 7809
rect 2593 7800 2605 7803
rect 2556 7772 2605 7800
rect 2556 7760 2562 7772
rect 2593 7769 2605 7772
rect 2639 7769 2651 7803
rect 2593 7763 2651 7769
rect 2685 7803 2743 7809
rect 2685 7769 2697 7803
rect 2731 7800 2743 7803
rect 4264 7800 4292 7828
rect 4540 7800 4568 7831
rect 4890 7828 4896 7880
rect 4948 7828 4954 7880
rect 5258 7828 5264 7880
rect 5316 7828 5322 7880
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5408 7840 5549 7868
rect 5408 7828 5414 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 2731 7772 4568 7800
rect 2731 7769 2743 7772
rect 2685 7763 2743 7769
rect 4982 7760 4988 7812
rect 5040 7760 5046 7812
rect 5123 7803 5181 7809
rect 5123 7769 5135 7803
rect 5169 7800 5181 7803
rect 5169 7772 5396 7800
rect 5169 7769 5181 7772
rect 5123 7763 5181 7769
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 1728 7704 2053 7732
rect 1728 7692 1734 7704
rect 2041 7701 2053 7704
rect 2087 7701 2099 7735
rect 2041 7695 2099 7701
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 5368 7741 5396 7772
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5644 7800 5672 7831
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 7392 7868 7420 7896
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7392 7840 7573 7868
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 7834 7868 7840 7880
rect 7699 7840 7840 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 5500 7772 5672 7800
rect 5905 7803 5963 7809
rect 5500 7760 5506 7772
rect 5905 7769 5917 7803
rect 5951 7800 5963 7803
rect 6270 7800 6276 7812
rect 5951 7772 6276 7800
rect 5951 7769 5963 7772
rect 5905 7763 5963 7769
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 7576 7800 7604 7831
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 7944 7877 7972 7976
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8202 7868 8208 7880
rect 8159 7840 8208 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8128 7800 8156 7831
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8352 7840 8401 7868
rect 8352 7828 8358 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 7024 7772 7420 7800
rect 7576 7772 8156 7800
rect 7024 7744 7052 7772
rect 4341 7735 4399 7741
rect 4341 7732 4353 7735
rect 4304 7704 4353 7732
rect 4304 7692 4310 7704
rect 4341 7701 4353 7704
rect 4387 7701 4399 7735
rect 4341 7695 4399 7701
rect 5353 7735 5411 7741
rect 5353 7701 5365 7735
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 7006 7692 7012 7744
rect 7064 7692 7070 7744
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 7392 7732 7420 7772
rect 7650 7732 7656 7744
rect 7392 7704 7656 7732
rect 7650 7692 7656 7704
rect 7708 7732 7714 7744
rect 8113 7735 8171 7741
rect 8113 7732 8125 7735
rect 7708 7704 8125 7732
rect 7708 7692 7714 7704
rect 8113 7701 8125 7704
rect 8159 7732 8171 7735
rect 8202 7732 8208 7744
rect 8159 7704 8208 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 8938 7732 8944 7744
rect 8619 7704 8944 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 1104 7642 9016 7664
rect 1104 7590 2599 7642
rect 2651 7590 2663 7642
rect 2715 7590 2727 7642
rect 2779 7590 2791 7642
rect 2843 7590 2855 7642
rect 2907 7590 4577 7642
rect 4629 7590 4641 7642
rect 4693 7590 4705 7642
rect 4757 7590 4769 7642
rect 4821 7590 4833 7642
rect 4885 7590 6555 7642
rect 6607 7590 6619 7642
rect 6671 7590 6683 7642
rect 6735 7590 6747 7642
rect 6799 7590 6811 7642
rect 6863 7590 8533 7642
rect 8585 7590 8597 7642
rect 8649 7590 8661 7642
rect 8713 7590 8725 7642
rect 8777 7590 8789 7642
rect 8841 7590 9016 7642
rect 1104 7568 9016 7590
rect 1854 7488 1860 7540
rect 1912 7488 1918 7540
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 2406 7528 2412 7540
rect 2271 7500 2412 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5258 7528 5264 7540
rect 4939 7500 5264 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 7190 7528 7196 7540
rect 6472 7500 7196 7528
rect 1670 7420 1676 7472
rect 1728 7469 1734 7472
rect 1728 7463 1777 7469
rect 1728 7429 1731 7463
rect 1765 7429 1777 7463
rect 1872 7460 1900 7488
rect 1949 7463 2007 7469
rect 1949 7460 1961 7463
rect 1872 7432 1961 7460
rect 1728 7423 1777 7429
rect 1949 7429 1961 7432
rect 1995 7429 2007 7463
rect 1949 7423 2007 7429
rect 4525 7463 4583 7469
rect 4525 7429 4537 7463
rect 4571 7460 4583 7463
rect 5460 7460 5488 7488
rect 4571 7432 5488 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 1728 7420 1734 7423
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1688 7364 1869 7392
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 1688 7324 1716 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 2041 7355 2099 7361
rect 4540 7364 4721 7392
rect 1544 7296 1716 7324
rect 1544 7284 1550 7296
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 2056 7324 2084 7355
rect 4540 7336 4568 7364
rect 4709 7361 4721 7364
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6472 7392 6500 7500
rect 7190 7488 7196 7500
rect 7248 7528 7254 7540
rect 7248 7500 7604 7528
rect 7248 7488 7254 7500
rect 6549 7463 6607 7469
rect 6549 7429 6561 7463
rect 6595 7460 6607 7463
rect 7576 7460 7604 7500
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 7834 7460 7840 7472
rect 6595 7432 7420 7460
rect 7576 7432 7840 7460
rect 6595 7429 6607 7432
rect 6549 7423 6607 7429
rect 6043 7364 6500 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 6914 7392 6920 7404
rect 6871 7364 6920 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7392 7401 7420 7432
rect 7834 7420 7840 7432
rect 7892 7460 7898 7472
rect 8021 7463 8079 7469
rect 8021 7460 8033 7463
rect 7892 7432 8033 7460
rect 7892 7420 7898 7432
rect 8021 7429 8033 7432
rect 8067 7429 8079 7463
rect 8021 7423 8079 7429
rect 7280 7395 7338 7401
rect 7280 7361 7292 7395
rect 7326 7361 7338 7395
rect 7280 7355 7338 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7367 7604 7395
rect 7515 7361 7527 7367
rect 7469 7355 7527 7361
rect 1820 7296 2084 7324
rect 1820 7284 1826 7296
rect 4522 7284 4528 7336
rect 4580 7284 4586 7336
rect 4982 7284 4988 7336
rect 5040 7324 5046 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 5040 7296 5273 7324
rect 5040 7284 5046 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 7300 7324 7328 7355
rect 7576 7336 7604 7367
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8478 7392 8484 7404
rect 8352 7364 8484 7392
rect 8352 7352 8358 7364
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 8570 7352 8576 7404
rect 8628 7352 8634 7404
rect 7300 7296 7512 7324
rect 5261 7287 5319 7293
rect 7484 7268 7512 7296
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 7466 7216 7472 7268
rect 7524 7216 7530 7268
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 8386 7188 8392 7200
rect 7055 7160 8392 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 1104 7098 9016 7120
rect 1104 7046 1939 7098
rect 1991 7046 2003 7098
rect 2055 7046 2067 7098
rect 2119 7046 2131 7098
rect 2183 7046 2195 7098
rect 2247 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 5895 7098
rect 5947 7046 5959 7098
rect 6011 7046 6023 7098
rect 6075 7046 6087 7098
rect 6139 7046 6151 7098
rect 6203 7046 7873 7098
rect 7925 7046 7937 7098
rect 7989 7046 8001 7098
rect 8053 7046 8065 7098
rect 8117 7046 8129 7098
rect 8181 7046 9016 7098
rect 1104 7024 9016 7046
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 4154 6984 4160 6996
rect 3467 6956 4160 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 4154 6944 4160 6956
rect 4212 6984 4218 6996
rect 4338 6984 4344 6996
rect 4212 6956 4344 6984
rect 4212 6944 4218 6956
rect 4338 6944 4344 6956
rect 4396 6984 4402 6996
rect 4525 6987 4583 6993
rect 4525 6984 4537 6987
rect 4396 6956 4537 6984
rect 4396 6944 4402 6956
rect 4525 6953 4537 6956
rect 4571 6953 4583 6987
rect 4525 6947 4583 6953
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 7098 6984 7104 6996
rect 5960 6956 7104 6984
rect 5960 6944 5966 6956
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 7282 6944 7288 6996
rect 7340 6944 7346 6996
rect 5442 6916 5448 6928
rect 5276 6888 5448 6916
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1949 6783 2007 6789
rect 1719 6752 1808 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 842 6604 848 6656
rect 900 6644 906 6656
rect 1780 6653 1808 6752
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2222 6780 2228 6792
rect 1995 6752 2228 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3252 6752 3985 6780
rect 2314 6672 2320 6724
rect 2372 6672 2378 6724
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 2501 6715 2559 6721
rect 2501 6712 2513 6715
rect 2464 6684 2513 6712
rect 2464 6672 2470 6684
rect 2501 6681 2513 6684
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 3252 6721 3280 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 5169 6783 5227 6789
rect 4304 6752 4752 6780
rect 4304 6740 4310 6752
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 3016 6684 3249 6712
rect 3016 6672 3022 6684
rect 3237 6681 3249 6684
rect 3283 6681 3295 6715
rect 3237 6675 3295 6681
rect 3528 6684 4016 6712
rect 1489 6647 1547 6653
rect 1489 6644 1501 6647
rect 900 6616 1501 6644
rect 900 6604 906 6616
rect 1489 6613 1501 6616
rect 1535 6613 1547 6647
rect 1489 6607 1547 6613
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6613 1823 6647
rect 1765 6607 1823 6613
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1912 6616 2145 6644
rect 1912 6604 1918 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 3442 6647 3500 6653
rect 3442 6613 3454 6647
rect 3488 6644 3500 6647
rect 3528 6644 3556 6684
rect 3488 6616 3556 6644
rect 3488 6613 3500 6616
rect 3442 6607 3500 6613
rect 3602 6604 3608 6656
rect 3660 6604 3666 6656
rect 3786 6604 3792 6656
rect 3844 6604 3850 6656
rect 3988 6644 4016 6684
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 4724 6721 4752 6752
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5276 6780 5304 6888
rect 5442 6876 5448 6888
rect 5500 6916 5506 6928
rect 5721 6919 5779 6925
rect 5721 6916 5733 6919
rect 5500 6888 5733 6916
rect 5500 6876 5506 6888
rect 5721 6885 5733 6888
rect 5767 6885 5779 6919
rect 5721 6879 5779 6885
rect 6454 6876 6460 6928
rect 6512 6876 6518 6928
rect 6914 6876 6920 6928
rect 6972 6916 6978 6928
rect 7745 6919 7803 6925
rect 7745 6916 7757 6919
rect 6972 6888 7757 6916
rect 6972 6876 6978 6888
rect 7745 6885 7757 6888
rect 7791 6885 7803 6919
rect 7745 6879 7803 6885
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 6472 6848 6500 6876
rect 5399 6820 6500 6848
rect 7668 6820 8340 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 6362 6780 6368 6792
rect 5215 6752 6368 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 6362 6740 6368 6752
rect 6420 6780 6426 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 6420 6752 6469 6780
rect 6420 6740 6426 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 6914 6783 6972 6789
rect 6914 6780 6926 6783
rect 6687 6752 6926 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 6914 6749 6926 6752
rect 6960 6780 6972 6783
rect 7190 6780 7196 6792
rect 6960 6752 7196 6780
rect 6960 6749 6972 6752
rect 6914 6743 6972 6749
rect 4493 6715 4551 6721
rect 4493 6712 4505 6715
rect 4120 6684 4505 6712
rect 4120 6672 4126 6684
rect 4493 6681 4505 6684
rect 4539 6681 4551 6715
rect 4493 6675 4551 6681
rect 4709 6715 4767 6721
rect 4709 6681 4721 6715
rect 4755 6681 4767 6715
rect 4709 6675 4767 6681
rect 4985 6715 5043 6721
rect 4985 6681 4997 6715
rect 5031 6712 5043 6715
rect 5074 6712 5080 6724
rect 5031 6684 5080 6712
rect 5031 6681 5043 6684
rect 4985 6675 5043 6681
rect 5074 6672 5080 6684
rect 5132 6712 5138 6724
rect 5350 6712 5356 6724
rect 5132 6684 5356 6712
rect 5132 6672 5138 6684
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 5810 6712 5816 6724
rect 5491 6684 5816 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5810 6672 5816 6684
rect 5868 6712 5874 6724
rect 6656 6712 6684 6743
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7668 6780 7696 6820
rect 7524 6752 7696 6780
rect 7524 6740 7530 6752
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8312 6789 8340 6820
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 8168 6752 8217 6780
rect 8168 6740 8174 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 7098 6712 7104 6724
rect 5868 6684 6684 6712
rect 6748 6684 7104 6712
rect 5868 6672 5874 6684
rect 4246 6644 4252 6656
rect 3988 6616 4252 6644
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 4338 6604 4344 6656
rect 4396 6604 4402 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 5718 6644 5724 6656
rect 4672 6616 5724 6644
rect 4672 6604 4678 6616
rect 5718 6604 5724 6616
rect 5776 6644 5782 6656
rect 5902 6644 5908 6656
rect 5776 6616 5908 6644
rect 5776 6604 5782 6616
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 6748 6653 6776 6684
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 8496 6712 8524 6743
rect 7616 6684 8524 6712
rect 8665 6715 8723 6721
rect 7616 6672 7622 6684
rect 8665 6681 8677 6715
rect 8711 6712 8723 6715
rect 8938 6712 8944 6724
rect 8711 6684 8944 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 8938 6672 8944 6684
rect 8996 6712 9002 6724
rect 9122 6712 9128 6724
rect 8996 6684 9128 6712
rect 8996 6672 9002 6684
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 6052 6616 6377 6644
rect 6052 6604 6058 6616
rect 6365 6613 6377 6616
rect 6411 6613 6423 6647
rect 6365 6607 6423 6613
rect 6733 6647 6791 6653
rect 6733 6613 6745 6647
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 6914 6604 6920 6656
rect 6972 6604 6978 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 8478 6644 8484 6656
rect 7064 6616 8484 6644
rect 7064 6604 7070 6616
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 1104 6554 9016 6576
rect 1104 6502 2599 6554
rect 2651 6502 2663 6554
rect 2715 6502 2727 6554
rect 2779 6502 2791 6554
rect 2843 6502 2855 6554
rect 2907 6502 4577 6554
rect 4629 6502 4641 6554
rect 4693 6502 4705 6554
rect 4757 6502 4769 6554
rect 4821 6502 4833 6554
rect 4885 6502 6555 6554
rect 6607 6502 6619 6554
rect 6671 6502 6683 6554
rect 6735 6502 6747 6554
rect 6799 6502 6811 6554
rect 6863 6502 8533 6554
rect 8585 6502 8597 6554
rect 8649 6502 8661 6554
rect 8713 6502 8725 6554
rect 8777 6502 8789 6554
rect 8841 6502 9016 6554
rect 1104 6480 9016 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 2590 6440 2596 6452
rect 2372 6412 2596 6440
rect 2372 6400 2378 6412
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2746 6412 2973 6440
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 1765 6375 1823 6381
rect 1765 6372 1777 6375
rect 1452 6344 1777 6372
rect 1452 6332 1458 6344
rect 1765 6341 1777 6344
rect 1811 6341 1823 6375
rect 1765 6335 1823 6341
rect 1949 6375 2007 6381
rect 1949 6341 1961 6375
rect 1995 6372 2007 6375
rect 2746 6372 2774 6412
rect 2961 6409 2973 6412
rect 3007 6440 3019 6443
rect 4062 6440 4068 6452
rect 3007 6412 4068 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 6089 6443 6147 6449
rect 6089 6409 6101 6443
rect 6135 6440 6147 6443
rect 6270 6440 6276 6452
rect 6135 6412 6276 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6270 6400 6276 6412
rect 6328 6440 6334 6452
rect 6638 6440 6644 6452
rect 6328 6412 6644 6440
rect 6328 6400 6334 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8478 6440 8484 6452
rect 8168 6412 8484 6440
rect 8168 6400 8174 6412
rect 8478 6400 8484 6412
rect 8536 6440 8542 6452
rect 9030 6440 9036 6452
rect 8536 6412 9036 6440
rect 8536 6400 8542 6412
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 3053 6375 3111 6381
rect 3053 6372 3065 6375
rect 1995 6344 2774 6372
rect 2884 6344 3065 6372
rect 1995 6341 2007 6344
rect 1949 6335 2007 6341
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2332 6313 2360 6344
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 2188 6276 2237 6304
rect 2188 6264 2194 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 2240 6168 2268 6267
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 2884 6304 2912 6344
rect 3053 6341 3065 6344
rect 3099 6341 3111 6375
rect 3053 6335 3111 6341
rect 3142 6332 3148 6384
rect 3200 6372 3206 6384
rect 4982 6372 4988 6384
rect 3200 6344 4988 6372
rect 3200 6332 3206 6344
rect 2832 6276 2912 6304
rect 2832 6264 2838 6276
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 3016 6276 3249 6304
rect 3016 6264 3022 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 4338 6304 4344 6316
rect 4111 6276 4344 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4908 6313 4936 6344
rect 4982 6332 4988 6344
rect 5040 6332 5046 6384
rect 7098 6372 7104 6384
rect 5276 6344 7104 6372
rect 5276 6313 5304 6344
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 2516 6236 2544 6264
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2516 6208 2605 6236
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 2731 6208 3433 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 3421 6205 3433 6208
rect 3467 6236 3479 6239
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3467 6208 3525 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4246 6236 4252 6248
rect 4019 6208 4252 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 2498 6168 2504 6180
rect 2240 6140 2504 6168
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 2608 6168 2636 6199
rect 2608 6140 2728 6168
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6100 1639 6103
rect 1670 6100 1676 6112
rect 1627 6072 1676 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 1820 6072 2053 6100
rect 1820 6060 1826 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2700 6100 2728 6140
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3712 6168 3740 6199
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 4448 6236 4476 6267
rect 4356 6208 4476 6236
rect 4908 6236 4936 6267
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5408 6276 5549 6304
rect 5408 6264 5414 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 5951 6276 6469 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6914 6304 6920 6316
rect 6604 6276 6920 6304
rect 6604 6264 6610 6276
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6304 7343 6307
rect 8128 6304 8156 6400
rect 7331 6276 8156 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 5626 6236 5632 6248
rect 4908 6208 5632 6236
rect 3108 6140 3740 6168
rect 3108 6128 3114 6140
rect 2774 6100 2780 6112
rect 2700 6072 2780 6100
rect 2041 6063 2099 6069
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 4356 6100 4384 6208
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6328 6208 6653 6236
rect 6328 6196 6334 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 5491 6140 5672 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 4890 6100 4896 6112
rect 3568 6072 4896 6100
rect 3568 6060 3574 6072
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 5040 6072 5089 6100
rect 5040 6060 5046 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5644 6100 5672 6140
rect 6362 6128 6368 6180
rect 6420 6168 6426 6180
rect 8036 6168 8064 6199
rect 6420 6140 8064 6168
rect 6420 6128 6426 6140
rect 7006 6100 7012 6112
rect 5644 6072 7012 6100
rect 5077 6063 5135 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7101 6103 7159 6109
rect 7101 6069 7113 6103
rect 7147 6100 7159 6103
rect 7650 6100 7656 6112
rect 7147 6072 7656 6100
rect 7147 6069 7159 6072
rect 7101 6063 7159 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 7742 6060 7748 6112
rect 7800 6060 7806 6112
rect 1104 6010 9016 6032
rect 1104 5958 1939 6010
rect 1991 5958 2003 6010
rect 2055 5958 2067 6010
rect 2119 5958 2131 6010
rect 2183 5958 2195 6010
rect 2247 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 5895 6010
rect 5947 5958 5959 6010
rect 6011 5958 6023 6010
rect 6075 5958 6087 6010
rect 6139 5958 6151 6010
rect 6203 5958 7873 6010
rect 7925 5958 7937 6010
rect 7989 5958 8001 6010
rect 8053 5958 8065 6010
rect 8117 5958 8129 6010
rect 8181 5958 9016 6010
rect 1104 5936 9016 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 3510 5896 3516 5908
rect 1627 5868 3516 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3660 5868 3893 5896
rect 3660 5856 3666 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 5166 5896 5172 5908
rect 4304 5868 5172 5896
rect 4304 5856 4310 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5902 5896 5908 5908
rect 5776 5868 5908 5896
rect 5776 5856 5782 5868
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 7432 5868 8493 5896
rect 7432 5856 7438 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 2464 5800 2636 5828
rect 2464 5788 2470 5800
rect 1670 5720 1676 5772
rect 1728 5720 1734 5772
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2501 5763 2559 5769
rect 2501 5760 2513 5763
rect 1912 5732 2084 5760
rect 1912 5720 1918 5732
rect 842 5652 848 5704
rect 900 5692 906 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 900 5664 1409 5692
rect 900 5652 906 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 2056 5701 2084 5732
rect 2148 5732 2513 5760
rect 2148 5701 2176 5732
rect 2501 5729 2513 5732
rect 2547 5729 2559 5763
rect 2501 5723 2559 5729
rect 2608 5760 2636 5800
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 7926 5828 7932 5840
rect 5868 5800 7932 5828
rect 5868 5788 5874 5800
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 8938 5828 8944 5840
rect 8220 5800 8944 5828
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 2608 5732 4261 5760
rect 2041 5695 2099 5701
rect 1544 5664 1992 5692
rect 1544 5652 1550 5664
rect 1964 5636 1992 5664
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 2406 5652 2412 5704
rect 2464 5652 2470 5704
rect 2608 5701 2636 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4338 5720 4344 5772
rect 4396 5720 4402 5772
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 5307 5732 7021 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 7009 5729 7021 5732
rect 7055 5760 7067 5763
rect 7466 5760 7472 5772
rect 7055 5732 7472 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8220 5769 8248 5800
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 8113 5763 8171 5769
rect 8113 5760 8125 5763
rect 7800 5732 8125 5760
rect 7800 5720 7806 5732
rect 8113 5729 8125 5732
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5729 8447 5763
rect 8389 5723 8447 5729
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 1762 5584 1768 5636
rect 1820 5633 1826 5636
rect 1820 5627 1869 5633
rect 1820 5593 1823 5627
rect 1857 5593 1869 5627
rect 1820 5587 1869 5593
rect 1820 5584 1826 5587
rect 1946 5584 1952 5636
rect 2004 5624 2010 5636
rect 3142 5624 3148 5636
rect 2004 5596 3148 5624
rect 2004 5584 2010 5596
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2682 5556 2688 5568
rect 2464 5528 2688 5556
rect 2464 5516 2470 5528
rect 2682 5516 2688 5528
rect 2740 5556 2746 5568
rect 3252 5556 3280 5655
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 4430 5652 4436 5704
rect 4488 5652 4494 5704
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5350 5692 5356 5704
rect 4847 5664 5356 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 4632 5624 4660 5655
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 6362 5692 6368 5704
rect 5675 5664 6368 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 7098 5692 7104 5704
rect 6687 5664 7104 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 4304 5596 4660 5624
rect 4304 5584 4310 5596
rect 4890 5584 4896 5636
rect 4948 5624 4954 5636
rect 4985 5627 5043 5633
rect 4985 5624 4997 5627
rect 4948 5596 4997 5624
rect 4948 5584 4954 5596
rect 4985 5593 4997 5596
rect 5031 5593 5043 5627
rect 4985 5587 5043 5593
rect 5442 5584 5448 5636
rect 5500 5584 5506 5636
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 5902 5624 5908 5636
rect 5592 5596 5908 5624
rect 5592 5584 5598 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 6089 5627 6147 5633
rect 6089 5593 6101 5627
rect 6135 5624 6147 5627
rect 6656 5624 6684 5655
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7432 5664 7665 5692
rect 7432 5652 7438 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8018 5652 8024 5704
rect 8076 5652 8082 5704
rect 8404 5692 8432 5723
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8404 5664 8493 5692
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 6135 5596 6684 5624
rect 6135 5593 6147 5596
rect 6089 5587 6147 5593
rect 6914 5584 6920 5636
rect 6972 5584 6978 5636
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7944 5624 7972 5652
rect 7524 5596 7972 5624
rect 7524 5584 7530 5596
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 8680 5624 8708 5655
rect 8444 5596 8708 5624
rect 8444 5584 8450 5596
rect 2740 5528 3280 5556
rect 3329 5559 3387 5565
rect 2740 5516 2746 5528
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3418 5556 3424 5568
rect 3375 5528 3424 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 5074 5516 5080 5568
rect 5132 5516 5138 5568
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 5994 5556 6000 5568
rect 5767 5528 6000 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6178 5516 6184 5568
rect 6236 5556 6242 5568
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 6236 5528 6377 5556
rect 6236 5516 6242 5528
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 7190 5516 7196 5568
rect 7248 5516 7254 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8478 5556 8484 5568
rect 8260 5528 8484 5556
rect 8260 5516 8266 5528
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 1104 5466 9016 5488
rect 1104 5414 2599 5466
rect 2651 5414 2663 5466
rect 2715 5414 2727 5466
rect 2779 5414 2791 5466
rect 2843 5414 2855 5466
rect 2907 5414 4577 5466
rect 4629 5414 4641 5466
rect 4693 5414 4705 5466
rect 4757 5414 4769 5466
rect 4821 5414 4833 5466
rect 4885 5414 6555 5466
rect 6607 5414 6619 5466
rect 6671 5414 6683 5466
rect 6735 5414 6747 5466
rect 6799 5414 6811 5466
rect 6863 5414 8533 5466
rect 8585 5414 8597 5466
rect 8649 5414 8661 5466
rect 8713 5414 8725 5466
rect 8777 5414 8789 5466
rect 8841 5414 9016 5466
rect 1104 5392 9016 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2406 5352 2412 5364
rect 1995 5324 2412 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 4246 5312 4252 5364
rect 4304 5312 4310 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5684 5324 5856 5352
rect 5684 5312 5690 5324
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 3786 5284 3792 5296
rect 992 5256 1808 5284
rect 992 5244 998 5256
rect 1780 5225 1808 5256
rect 3344 5256 3792 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2314 5216 2320 5228
rect 2271 5188 2320 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 1688 5148 1716 5179
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 3344 5225 3372 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 4798 5244 4804 5296
rect 4856 5284 4862 5296
rect 4856 5256 5580 5284
rect 4856 5244 4862 5256
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3418 5176 3424 5228
rect 3476 5176 3482 5228
rect 3602 5176 3608 5228
rect 3660 5176 3666 5228
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4338 5216 4344 5228
rect 4203 5188 4344 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4614 5216 4620 5228
rect 4571 5188 4620 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 5074 5216 5080 5228
rect 4816 5188 5080 5216
rect 1688 5120 2084 5148
rect 2056 5089 2084 5120
rect 2498 5108 2504 5160
rect 2556 5148 2562 5160
rect 4433 5151 4491 5157
rect 4433 5148 4445 5151
rect 2556 5120 4445 5148
rect 2556 5108 2562 5120
rect 4433 5117 4445 5120
rect 4479 5148 4491 5151
rect 4816 5148 4844 5188
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5215 5188 5457 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 4479 5120 4844 5148
rect 4893 5151 4951 5157
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 4893 5117 4905 5151
rect 4939 5148 4951 5151
rect 4982 5148 4988 5160
rect 4939 5120 4988 5148
rect 4939 5117 4951 5120
rect 4893 5111 4951 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5552 5148 5580 5256
rect 5626 5177 5632 5229
rect 5684 5177 5690 5229
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 5828 5225 5856 5324
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6144 5324 6377 5352
rect 6144 5312 6150 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 5994 5293 6000 5296
rect 5951 5287 6000 5293
rect 5951 5253 5963 5287
rect 5997 5253 6000 5287
rect 5951 5247 6000 5253
rect 5994 5244 6000 5247
rect 6052 5244 6058 5296
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5216 6147 5219
rect 6178 5216 6184 5228
rect 6135 5188 6184 5216
rect 6135 5185 6147 5188
rect 6089 5179 6147 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6730 5216 6736 5228
rect 6595 5188 6736 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 6932 5188 7297 5216
rect 6822 5148 6828 5160
rect 5552 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 6932 5092 6960 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7285 5179 7343 5185
rect 7392 5188 7665 5216
rect 7392 5148 7420 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7300 5120 7420 5148
rect 7300 5092 7328 5120
rect 2041 5083 2099 5089
rect 2041 5049 2053 5083
rect 2087 5049 2099 5083
rect 2041 5043 2099 5049
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6914 5080 6920 5092
rect 5500 5052 6920 5080
rect 5500 5040 5506 5052
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7282 5040 7288 5092
rect 7340 5040 7346 5092
rect 7374 5040 7380 5092
rect 7432 5040 7438 5092
rect 1486 4972 1492 5024
rect 1544 4972 1550 5024
rect 3142 4972 3148 5024
rect 3200 4972 3206 5024
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3752 4984 3985 5012
rect 3752 4972 3758 4984
rect 3973 4981 3985 4984
rect 4019 4981 4031 5015
rect 3973 4975 4031 4981
rect 5353 5015 5411 5021
rect 5353 4981 5365 5015
rect 5399 5012 5411 5015
rect 8386 5012 8392 5024
rect 5399 4984 8392 5012
rect 5399 4981 5411 4984
rect 5353 4975 5411 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 1104 4922 9016 4944
rect 1104 4870 1939 4922
rect 1991 4870 2003 4922
rect 2055 4870 2067 4922
rect 2119 4870 2131 4922
rect 2183 4870 2195 4922
rect 2247 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 5895 4922
rect 5947 4870 5959 4922
rect 6011 4870 6023 4922
rect 6075 4870 6087 4922
rect 6139 4870 6151 4922
rect 6203 4870 7873 4922
rect 7925 4870 7937 4922
rect 7989 4870 8001 4922
rect 8053 4870 8065 4922
rect 8117 4870 8129 4922
rect 8181 4870 9016 4922
rect 1104 4848 9016 4870
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4614 4808 4620 4820
rect 4212 4780 4620 4808
rect 4212 4768 4218 4780
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 8352 4780 8493 4808
rect 8352 4768 8358 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 2958 4740 2964 4752
rect 2608 4712 2964 4740
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4672 2283 4675
rect 2498 4672 2504 4684
rect 2271 4644 2504 4672
rect 2271 4641 2283 4644
rect 2225 4635 2283 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 2608 4681 2636 4712
rect 2958 4700 2964 4712
rect 3016 4740 3022 4752
rect 4798 4740 4804 4752
rect 3016 4712 4804 4740
rect 3016 4700 3022 4712
rect 4798 4700 4804 4712
rect 4856 4700 4862 4752
rect 5258 4700 5264 4752
rect 5316 4700 5322 4752
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 5736 4712 7481 4740
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4641 2651 4675
rect 2593 4635 2651 4641
rect 4246 4632 4252 4684
rect 4304 4632 4310 4684
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5736 4681 5764 4712
rect 7469 4709 7481 4712
rect 7515 4709 7527 4743
rect 7469 4703 7527 4709
rect 5721 4675 5779 4681
rect 5721 4672 5733 4675
rect 5224 4644 5733 4672
rect 5224 4632 5230 4644
rect 5721 4641 5733 4644
rect 5767 4641 5779 4675
rect 5721 4635 5779 4641
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 5868 4644 6040 4672
rect 5868 4632 5874 4644
rect 1394 4564 1400 4616
rect 1452 4604 1458 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1452 4576 1777 4604
rect 1452 4564 1458 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2685 4607 2743 4613
rect 2363 4576 2397 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2958 4604 2964 4616
rect 2731 4576 2964 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 1949 4539 2007 4545
rect 1949 4505 1961 4539
rect 1995 4536 2007 4539
rect 2332 4536 2360 4567
rect 2958 4564 2964 4576
rect 3016 4604 3022 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3016 4576 3801 4604
rect 3016 4564 3022 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 6012 4613 6040 4644
rect 6270 4632 6276 4684
rect 6328 4632 6334 4684
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7285 4675 7343 4681
rect 7285 4672 7297 4675
rect 7248 4644 7297 4672
rect 7248 4632 7254 4644
rect 7285 4641 7297 4644
rect 7331 4641 7343 4675
rect 7285 4635 7343 4641
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7708 4644 8033 4672
rect 7708 4632 7714 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 6288 4604 6316 4632
rect 7742 4604 7748 4616
rect 6288 4576 7748 4604
rect 5997 4567 6055 4573
rect 7742 4564 7748 4576
rect 7800 4604 7806 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7800 4576 7941 4604
rect 7800 4564 7806 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 2406 4536 2412 4548
rect 1995 4508 2412 4536
rect 1995 4505 2007 4508
rect 1949 4499 2007 4505
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 3602 4496 3608 4548
rect 3660 4536 3666 4548
rect 4890 4536 4896 4548
rect 3660 4508 4896 4536
rect 3660 4496 3666 4508
rect 4890 4496 4896 4508
rect 4948 4536 4954 4548
rect 4948 4508 5028 4536
rect 4948 4496 4954 4508
rect 1578 4428 1584 4480
rect 1636 4428 1642 4480
rect 2038 4428 2044 4480
rect 2096 4428 2102 4480
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 3844 4440 3985 4468
rect 3844 4428 3850 4440
rect 3973 4437 3985 4440
rect 4019 4437 4031 4471
rect 5000 4468 5028 4508
rect 5074 4496 5080 4548
rect 5132 4536 5138 4548
rect 5813 4539 5871 4545
rect 5813 4536 5825 4539
rect 5132 4508 5825 4536
rect 5132 4496 5138 4508
rect 5813 4505 5825 4508
rect 5859 4505 5871 4539
rect 5813 4499 5871 4505
rect 5718 4468 5724 4480
rect 5000 4440 5724 4468
rect 3973 4431 4031 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 1104 4378 9016 4400
rect 1104 4326 2599 4378
rect 2651 4326 2663 4378
rect 2715 4326 2727 4378
rect 2779 4326 2791 4378
rect 2843 4326 2855 4378
rect 2907 4326 4577 4378
rect 4629 4326 4641 4378
rect 4693 4326 4705 4378
rect 4757 4326 4769 4378
rect 4821 4326 4833 4378
rect 4885 4326 6555 4378
rect 6607 4326 6619 4378
rect 6671 4326 6683 4378
rect 6735 4326 6747 4378
rect 6799 4326 6811 4378
rect 6863 4326 8533 4378
rect 8585 4326 8597 4378
rect 8649 4326 8661 4378
rect 8713 4326 8725 4378
rect 8777 4326 8789 4378
rect 8841 4326 9016 4378
rect 1104 4304 9016 4326
rect 2038 4224 2044 4276
rect 2096 4224 2102 4276
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 2314 4264 2320 4276
rect 2271 4236 2320 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2885 4267 2943 4273
rect 2885 4264 2897 4267
rect 2464 4236 2897 4264
rect 2464 4224 2470 4236
rect 2885 4233 2897 4236
rect 2931 4233 2943 4267
rect 2885 4227 2943 4233
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3292 4236 4216 4264
rect 3292 4224 3298 4236
rect 1739 4199 1797 4205
rect 1739 4165 1751 4199
rect 1785 4196 1797 4199
rect 2056 4196 2084 4224
rect 1785 4168 2084 4196
rect 2685 4199 2743 4205
rect 1785 4165 1797 4168
rect 1739 4159 1797 4165
rect 2685 4165 2697 4199
rect 2731 4165 2743 4199
rect 2685 4159 2743 4165
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 1946 4088 1952 4140
rect 2004 4088 2010 4140
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 2056 3992 2084 4091
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2700 4128 2728 4159
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 3602 4196 3608 4208
rect 2832 4168 3608 4196
rect 2832 4156 2838 4168
rect 3602 4156 3608 4168
rect 3660 4156 3666 4208
rect 4188 4196 4216 4236
rect 4246 4224 4252 4276
rect 4304 4224 4310 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4488 4236 4813 4264
rect 4488 4224 4494 4236
rect 4801 4233 4813 4236
rect 4847 4233 4859 4267
rect 4801 4227 4859 4233
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 5684 4236 6377 4264
rect 5684 4224 5690 4236
rect 6365 4233 6377 4236
rect 6411 4233 6423 4267
rect 6365 4227 6423 4233
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7098 4264 7104 4276
rect 7055 4236 7104 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7558 4224 7564 4276
rect 7616 4224 7622 4276
rect 5166 4196 5172 4208
rect 4188 4168 4568 4196
rect 3050 4128 3056 4140
rect 2556 4100 3056 4128
rect 2556 4088 2562 4100
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 4065 4131 4123 4137
rect 3528 4100 3924 4128
rect 1820 3964 2084 3992
rect 3053 3995 3111 4001
rect 1820 3952 1826 3964
rect 3053 3961 3065 3995
rect 3099 3992 3111 3995
rect 3528 3992 3556 4100
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3660 4032 3801 4060
rect 3660 4020 3666 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 3896 4060 3924 4100
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4430 4128 4436 4140
rect 4111 4100 4436 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4338 4060 4344 4072
rect 3896 4032 4344 4060
rect 3789 4023 3847 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 4540 4060 4568 4168
rect 4724 4168 5172 4196
rect 4724 4137 4752 4168
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 7190 4196 7196 4208
rect 6779 4168 7196 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4097 4767 4131
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 4709 4091 4767 4097
rect 4816 4100 5089 4128
rect 4816 4060 4844 4100
rect 5077 4097 5089 4100
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5350 4128 5356 4140
rect 5307 4100 5356 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 4540 4032 4844 4060
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 3099 3964 3556 3992
rect 3881 3995 3939 4001
rect 3099 3961 3111 3964
rect 3053 3955 3111 3961
rect 3881 3961 3893 3995
rect 3927 3992 3939 3995
rect 5000 3992 5028 4023
rect 5166 4020 5172 4072
rect 5224 4020 5230 4072
rect 5736 4060 5764 4091
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5868 4100 5917 4128
rect 5868 4088 5874 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 6178 4088 6184 4140
rect 6236 4088 6242 4140
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6420 4100 6561 4128
rect 6420 4088 6426 4100
rect 6549 4097 6561 4100
rect 6595 4128 6607 4131
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6595 4100 6837 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 6270 4060 6276 4072
rect 5736 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 3927 3964 5028 3992
rect 5997 3995 6055 4001
rect 3927 3961 3939 3964
rect 3881 3955 3939 3961
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 6362 3992 6368 4004
rect 6043 3964 6368 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 6840 3992 6868 4091
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 7024 4060 7052 4091
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7432 4100 7757 4128
rect 7432 4088 7438 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 6972 4032 7052 4060
rect 6972 4020 6978 4032
rect 7098 4020 7104 4072
rect 7156 4020 7162 4072
rect 7650 4020 7656 4072
rect 7708 4020 7714 4072
rect 7944 3992 7972 4091
rect 8202 4088 8208 4140
rect 8260 4088 8266 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 6840 3964 7972 3992
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 8938 3992 8944 4004
rect 8619 3964 8944 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2372 3896 2881 3924
rect 2372 3884 2378 3896
rect 2869 3893 2881 3896
rect 2915 3924 2927 3927
rect 3142 3924 3148 3936
rect 2915 3896 3148 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3326 3884 3332 3936
rect 3384 3924 3390 3936
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3384 3896 3985 3924
rect 3384 3884 3390 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 3973 3887 4031 3893
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5592 3896 5825 3924
rect 5592 3884 5598 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 1104 3834 9016 3856
rect 1104 3782 1939 3834
rect 1991 3782 2003 3834
rect 2055 3782 2067 3834
rect 2119 3782 2131 3834
rect 2183 3782 2195 3834
rect 2247 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 5895 3834
rect 5947 3782 5959 3834
rect 6011 3782 6023 3834
rect 6075 3782 6087 3834
rect 6139 3782 6151 3834
rect 6203 3782 7873 3834
rect 7925 3782 7937 3834
rect 7989 3782 8001 3834
rect 8053 3782 8065 3834
rect 8117 3782 8129 3834
rect 8181 3782 9016 3834
rect 1104 3760 9016 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 1857 3723 1915 3729
rect 1857 3720 1869 3723
rect 1820 3692 1869 3720
rect 1820 3680 1826 3692
rect 1857 3689 1869 3692
rect 1903 3689 1915 3723
rect 1857 3683 1915 3689
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2406 3720 2412 3732
rect 2179 3692 2412 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2958 3720 2964 3732
rect 2823 3692 2964 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 4028 3692 4169 3720
rect 4028 3680 4034 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 4157 3683 4215 3689
rect 5258 3680 5264 3732
rect 5316 3680 5322 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 8478 3720 8484 3732
rect 5684 3692 8484 3720
rect 5684 3680 5690 3692
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 3145 3655 3203 3661
rect 1627 3624 1992 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 1964 3596 1992 3624
rect 3145 3621 3157 3655
rect 3191 3621 3203 3655
rect 3145 3615 3203 3621
rect 4341 3655 4399 3661
rect 4341 3621 4353 3655
rect 4387 3652 4399 3655
rect 6549 3655 6607 3661
rect 4387 3624 5120 3652
rect 4387 3621 4399 3624
rect 4341 3615 4399 3621
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 3160 3584 3188 3615
rect 3510 3584 3516 3596
rect 2004 3556 2268 3584
rect 3160 3556 3516 3584
rect 2004 3544 2010 3556
rect 1394 3476 1400 3528
rect 1452 3476 1458 3528
rect 1670 3476 1676 3528
rect 1728 3476 1734 3528
rect 1762 3476 1768 3528
rect 1820 3476 1826 3528
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 2240 3525 2268 3556
rect 3510 3544 3516 3556
rect 3568 3584 3574 3596
rect 4062 3584 4068 3596
rect 3568 3556 4068 3584
rect 3568 3544 3574 3556
rect 4062 3544 4068 3556
rect 4120 3584 4126 3596
rect 4801 3587 4859 3593
rect 4120 3556 4660 3584
rect 4120 3544 4126 3556
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 2271 3488 2421 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2409 3485 2421 3488
rect 2455 3516 2467 3519
rect 2869 3519 2927 3525
rect 2869 3516 2881 3519
rect 2455 3488 2881 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 2869 3485 2881 3488
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3292 3488 3341 3516
rect 3292 3476 3298 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3786 3516 3792 3528
rect 3651 3488 3792 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 4632 3525 4660 3556
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 4982 3584 4988 3596
rect 4847 3556 4988 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 4908 3525 4936 3556
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 5092 3584 5120 3624
rect 5276 3624 5948 3652
rect 5276 3596 5304 3624
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 5092 3556 5181 3584
rect 5169 3553 5181 3556
rect 5215 3553 5227 3587
rect 5169 3547 5227 3553
rect 5258 3544 5264 3596
rect 5316 3544 5322 3596
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5920 3593 5948 3624
rect 6549 3621 6561 3655
rect 6595 3652 6607 3655
rect 6914 3652 6920 3664
rect 6595 3624 6920 3652
rect 6595 3621 6607 3624
rect 6549 3615 6607 3621
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7282 3612 7288 3664
rect 7340 3652 7346 3664
rect 8202 3652 8208 3664
rect 7340 3624 8208 3652
rect 7340 3612 7346 3624
rect 8202 3612 8208 3624
rect 8260 3652 8266 3664
rect 8260 3624 8432 3652
rect 8260 3612 8266 3624
rect 5905 3587 5963 3593
rect 5408 3556 5856 3584
rect 5408 3544 5414 3556
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3516 4951 3519
rect 5537 3519 5595 3525
rect 4939 3488 4973 3516
rect 4939 3485 4951 3488
rect 4893 3479 4951 3485
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 2056 3448 2084 3476
rect 2593 3451 2651 3457
rect 2593 3448 2605 3451
rect 2056 3420 2605 3448
rect 2593 3417 2605 3420
rect 2639 3417 2651 3451
rect 2593 3411 2651 3417
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 3973 3451 4031 3457
rect 3973 3448 3985 3451
rect 3936 3420 3985 3448
rect 3936 3408 3942 3420
rect 3973 3417 3985 3420
rect 4019 3417 4031 3451
rect 3973 3411 4031 3417
rect 4154 3408 4160 3460
rect 4212 3457 4218 3460
rect 4212 3451 4231 3457
rect 4219 3417 4231 3451
rect 4212 3411 4231 3417
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3417 4491 3451
rect 4433 3411 4491 3417
rect 4212 3408 4218 3411
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2774 3380 2780 3392
rect 2556 3352 2780 3380
rect 2556 3340 2562 3352
rect 2774 3340 2780 3352
rect 2832 3340 2838 3392
rect 2958 3340 2964 3392
rect 3016 3340 3022 3392
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3108 3352 3433 3380
rect 3108 3340 3114 3352
rect 3421 3349 3433 3352
rect 3467 3380 3479 3383
rect 3602 3380 3608 3392
rect 3467 3352 3608 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3602 3340 3608 3352
rect 3660 3380 3666 3392
rect 4338 3380 4344 3392
rect 3660 3352 4344 3380
rect 3660 3340 3666 3352
rect 4338 3340 4344 3352
rect 4396 3380 4402 3392
rect 4448 3380 4476 3411
rect 4522 3408 4528 3460
rect 4580 3448 4586 3460
rect 5552 3448 5580 3479
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 5828 3516 5856 3556
rect 5905 3553 5917 3587
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 8404 3593 8432 3624
rect 8389 3587 8447 3593
rect 7800 3556 7972 3584
rect 7800 3544 7806 3556
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 5828 3488 6193 3516
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 7006 3476 7012 3528
rect 7064 3476 7070 3528
rect 7190 3476 7196 3528
rect 7248 3476 7254 3528
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 4580 3420 5580 3448
rect 4580 3408 4586 3420
rect 4396 3352 4476 3380
rect 4396 3340 4402 3352
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 5445 3383 5503 3389
rect 5445 3380 5457 3383
rect 5132 3352 5457 3380
rect 5132 3340 5138 3352
rect 5445 3349 5457 3352
rect 5491 3349 5503 3383
rect 5445 3343 5503 3349
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 5629 3383 5687 3389
rect 5629 3380 5641 3383
rect 5592 3352 5641 3380
rect 5592 3340 5598 3352
rect 5629 3349 5641 3352
rect 5675 3349 5687 3383
rect 5736 3380 5764 3476
rect 6089 3451 6147 3457
rect 6089 3417 6101 3451
rect 6135 3448 6147 3451
rect 6362 3448 6368 3460
rect 6135 3420 6368 3448
rect 6135 3417 6147 3420
rect 6089 3411 6147 3417
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 7300 3448 7328 3479
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7944 3516 7972 3556
rect 8389 3553 8401 3587
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 8030 3519 8088 3525
rect 8030 3516 8042 3519
rect 7944 3488 8042 3516
rect 7837 3479 7895 3485
rect 8030 3485 8042 3488
rect 8076 3485 8088 3519
rect 8030 3479 8088 3485
rect 7742 3448 7748 3460
rect 6748 3420 7748 3448
rect 6748 3380 6776 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 7852 3448 7880 3479
rect 8386 3448 8392 3460
rect 7852 3420 8392 3448
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 5736 3352 6776 3380
rect 5629 3343 5687 3349
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 8110 3380 8116 3392
rect 6880 3352 8116 3380
rect 6880 3340 6886 3352
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 1104 3290 9016 3312
rect 1104 3238 2599 3290
rect 2651 3238 2663 3290
rect 2715 3238 2727 3290
rect 2779 3238 2791 3290
rect 2843 3238 2855 3290
rect 2907 3238 4577 3290
rect 4629 3238 4641 3290
rect 4693 3238 4705 3290
rect 4757 3238 4769 3290
rect 4821 3238 4833 3290
rect 4885 3238 6555 3290
rect 6607 3238 6619 3290
rect 6671 3238 6683 3290
rect 6735 3238 6747 3290
rect 6799 3238 6811 3290
rect 6863 3238 8533 3290
rect 8585 3238 8597 3290
rect 8649 3238 8661 3290
rect 8713 3238 8725 3290
rect 8777 3238 8789 3290
rect 8841 3238 9016 3290
rect 1104 3216 9016 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1912 3148 1961 3176
rect 1912 3136 1918 3148
rect 1949 3145 1961 3148
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 2056 3148 3372 3176
rect 2056 3120 2084 3148
rect 2038 3068 2044 3120
rect 2096 3068 2102 3120
rect 2257 3111 2315 3117
rect 2257 3077 2269 3111
rect 2303 3108 2315 3111
rect 2406 3108 2412 3120
rect 2303 3080 2412 3108
rect 2303 3077 2315 3080
rect 2257 3071 2315 3077
rect 2406 3068 2412 3080
rect 2464 3108 2470 3120
rect 2958 3108 2964 3120
rect 2464 3080 2728 3108
rect 2464 3068 2470 3080
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1762 3040 1768 3052
rect 1636 3012 1768 3040
rect 1636 3000 1642 3012
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2056 3040 2084 3068
rect 1912 3012 2084 3040
rect 1912 3000 1918 3012
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 1946 2972 1952 2984
rect 1719 2944 1952 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2608 2972 2636 3003
rect 2424 2944 2636 2972
rect 2700 2972 2728 3080
rect 2792 3080 2964 3108
rect 2792 3049 2820 3080
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 3344 3049 3372 3148
rect 3418 3136 3424 3188
rect 3476 3176 3482 3188
rect 3513 3179 3571 3185
rect 3513 3176 3525 3179
rect 3476 3148 3525 3176
rect 3476 3136 3482 3148
rect 3513 3145 3525 3148
rect 3559 3145 3571 3179
rect 3513 3139 3571 3145
rect 3602 3136 3608 3188
rect 3660 3136 3666 3188
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4430 3176 4436 3188
rect 4203 3148 4436 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 3620 3108 3648 3136
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 3620 3080 3801 3108
rect 3789 3077 3801 3080
rect 3835 3108 3847 3111
rect 3878 3108 3884 3120
rect 3835 3080 3884 3108
rect 3835 3077 3847 3080
rect 3789 3071 3847 3077
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 4062 3117 4068 3120
rect 4005 3111 4068 3117
rect 4005 3077 4017 3111
rect 4051 3077 4068 3111
rect 4005 3071 4068 3077
rect 4062 3068 4068 3071
rect 4120 3068 4126 3120
rect 4264 3049 4292 3148
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 5074 3136 5080 3188
rect 5132 3136 5138 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7374 3176 7380 3188
rect 6696 3148 7380 3176
rect 6696 3136 6702 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7834 3176 7840 3188
rect 7524 3148 7840 3176
rect 7524 3136 7530 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8294 3176 8300 3188
rect 8159 3148 8300 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 4985 3111 5043 3117
rect 4985 3077 4997 3111
rect 5031 3108 5043 3111
rect 5166 3108 5172 3120
rect 5031 3080 5172 3108
rect 5031 3077 5043 3080
rect 4985 3071 5043 3077
rect 5166 3068 5172 3080
rect 5224 3108 5230 3120
rect 8404 3108 8432 3139
rect 5224 3080 5488 3108
rect 5224 3068 5230 3080
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2915 3012 3157 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 3620 2972 3648 3003
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 5460 3049 5488 3080
rect 6196 3080 8432 3108
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4396 3012 4537 3040
rect 4396 3000 4402 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5534 3000 5540 3052
rect 5592 3000 5598 3052
rect 5626 3000 5632 3052
rect 5684 3000 5690 3052
rect 6196 3049 6224 3080
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 6638 3040 6644 3052
rect 6181 3003 6239 3009
rect 6380 3012 6644 3040
rect 2700 2944 3648 2972
rect 5644 2972 5672 3000
rect 6380 2972 6408 3012
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 6840 3012 7297 3040
rect 6840 2984 6868 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7742 3000 7748 3052
rect 7800 3000 7806 3052
rect 8110 3000 8116 3052
rect 8168 3000 8174 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8260 3012 8309 3040
rect 8260 3000 8266 3012
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 5644 2944 6408 2972
rect 6457 2975 6515 2981
rect 2424 2913 2452 2944
rect 6457 2941 6469 2975
rect 6503 2972 6515 2975
rect 6822 2972 6828 2984
rect 6503 2944 6828 2972
rect 6503 2941 6515 2944
rect 6457 2935 6515 2941
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7064 2944 7481 2972
rect 7064 2932 7070 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7834 2972 7840 2984
rect 7607 2944 7840 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 2409 2907 2467 2913
rect 2409 2904 2421 2907
rect 1688 2876 2421 2904
rect 1688 2848 1716 2876
rect 2409 2873 2421 2876
rect 2455 2873 2467 2907
rect 2409 2867 2467 2873
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 4154 2904 4160 2916
rect 2648 2876 4160 2904
rect 2648 2864 2654 2876
rect 4154 2864 4160 2876
rect 4212 2864 4218 2916
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 4430 2904 4436 2916
rect 4387 2876 4436 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 6917 2907 6975 2913
rect 6917 2873 6929 2907
rect 6963 2904 6975 2907
rect 6963 2876 7328 2904
rect 6963 2873 6975 2876
rect 6917 2867 6975 2873
rect 7300 2848 7328 2876
rect 1670 2796 1676 2848
rect 1728 2796 1734 2848
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2314 2836 2320 2848
rect 2271 2808 2320 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3510 2836 3516 2848
rect 3099 2808 3516 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3510 2796 3516 2808
rect 3568 2836 3574 2848
rect 3970 2836 3976 2848
rect 3568 2808 3976 2836
rect 3568 2796 3574 2808
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 5718 2796 5724 2848
rect 5776 2796 5782 2848
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6454 2836 6460 2848
rect 6043 2808 6460 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 7190 2836 7196 2848
rect 7147 2808 7196 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7282 2796 7288 2848
rect 7340 2796 7346 2848
rect 7484 2836 7512 2935
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 7742 2864 7748 2916
rect 7800 2904 7806 2916
rect 8588 2904 8616 3003
rect 7800 2876 8616 2904
rect 7800 2864 7806 2876
rect 8294 2836 8300 2848
rect 7484 2808 8300 2836
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 1104 2746 9016 2768
rect 1104 2694 1939 2746
rect 1991 2694 2003 2746
rect 2055 2694 2067 2746
rect 2119 2694 2131 2746
rect 2183 2694 2195 2746
rect 2247 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 5895 2746
rect 5947 2694 5959 2746
rect 6011 2694 6023 2746
rect 6075 2694 6087 2746
rect 6139 2694 6151 2746
rect 6203 2694 7873 2746
rect 7925 2694 7937 2746
rect 7989 2694 8001 2746
rect 8053 2694 8065 2746
rect 8117 2694 8129 2746
rect 8181 2694 9016 2746
rect 1104 2672 9016 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 1636 2604 1961 2632
rect 1636 2592 1642 2604
rect 1949 2601 1961 2604
rect 1995 2601 2007 2635
rect 1949 2595 2007 2601
rect 2222 2592 2228 2644
rect 2280 2632 2286 2644
rect 2406 2632 2412 2644
rect 2280 2604 2412 2632
rect 2280 2592 2286 2604
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 3050 2632 3056 2644
rect 2516 2604 3056 2632
rect 2406 2496 2412 2508
rect 1412 2468 2412 2496
rect 1412 2437 1440 2468
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 2222 2388 2228 2440
rect 2280 2388 2286 2440
rect 2516 2437 2544 2604
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3326 2592 3332 2644
rect 3384 2632 3390 2644
rect 4430 2632 4436 2644
rect 3384 2604 4436 2632
rect 3384 2592 3390 2604
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 6270 2632 6276 2644
rect 5592 2604 6276 2632
rect 5592 2592 5598 2604
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6362 2592 6368 2644
rect 6420 2592 6426 2644
rect 7006 2632 7012 2644
rect 6748 2604 7012 2632
rect 2590 2524 2596 2576
rect 2648 2524 2654 2576
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 5258 2564 5264 2576
rect 3191 2536 5264 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 5442 2524 5448 2576
rect 5500 2564 5506 2576
rect 6748 2573 6776 2604
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 7374 2632 7380 2644
rect 7239 2604 7380 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7558 2592 7564 2644
rect 7616 2632 7622 2644
rect 7653 2635 7711 2641
rect 7653 2632 7665 2635
rect 7616 2604 7665 2632
rect 7616 2592 7622 2604
rect 7653 2601 7665 2604
rect 7699 2601 7711 2635
rect 7653 2595 7711 2601
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 8444 2604 8493 2632
rect 8444 2592 8450 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 5500 2536 6745 2564
rect 5500 2524 5506 2536
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 7745 2567 7803 2573
rect 7745 2564 7757 2567
rect 6733 2527 6791 2533
rect 7024 2536 7757 2564
rect 5460 2496 5488 2524
rect 2700 2468 3188 2496
rect 2700 2437 2728 2468
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 2866 2428 2872 2440
rect 2823 2400 2872 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 1762 2360 1768 2372
rect 1596 2332 1768 2360
rect 1596 2301 1624 2332
rect 1762 2320 1768 2332
rect 1820 2360 1826 2372
rect 1949 2363 2007 2369
rect 1949 2360 1961 2363
rect 1820 2332 1961 2360
rect 1820 2320 1826 2332
rect 1949 2329 1961 2332
rect 1995 2329 2007 2363
rect 1949 2323 2007 2329
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 1854 2252 1860 2304
rect 1912 2252 1918 2304
rect 2133 2295 2191 2301
rect 2133 2261 2145 2295
rect 2179 2292 2191 2295
rect 2314 2292 2320 2304
rect 2179 2264 2320 2292
rect 2179 2261 2191 2264
rect 2133 2255 2191 2261
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 2961 2295 3019 2301
rect 2961 2261 2973 2295
rect 3007 2292 3019 2295
rect 3068 2292 3096 2391
rect 3160 2360 3188 2468
rect 3252 2468 5488 2496
rect 3252 2437 3280 2468
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 5592 2468 5856 2496
rect 5592 2456 5598 2468
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2428 3387 2431
rect 3418 2428 3424 2440
rect 3375 2400 3424 2428
rect 3375 2397 3387 2400
rect 3329 2391 3387 2397
rect 3344 2360 3372 2391
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 3510 2388 3516 2440
rect 3568 2388 3574 2440
rect 3602 2388 3608 2440
rect 3660 2388 3666 2440
rect 3694 2388 3700 2440
rect 3752 2428 3758 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3752 2400 4077 2428
rect 3752 2388 3758 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 5445 2431 5503 2437
rect 4212 2400 5396 2428
rect 4212 2388 4218 2400
rect 3160 2332 3372 2360
rect 4430 2320 4436 2372
rect 4488 2320 4494 2372
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5166 2360 5172 2372
rect 5123 2332 5172 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5166 2320 5172 2332
rect 5224 2320 5230 2372
rect 5368 2360 5396 2400
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5718 2428 5724 2440
rect 5491 2400 5724 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5828 2437 5856 2468
rect 6012 2468 6837 2496
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 6012 2369 6040 2468
rect 6825 2465 6837 2468
rect 6871 2496 6883 2499
rect 7024 2496 7052 2536
rect 7745 2533 7757 2536
rect 7791 2533 7803 2567
rect 7745 2527 7803 2533
rect 6871 2468 7052 2496
rect 6871 2465 6883 2468
rect 6825 2459 6883 2465
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 7524 2468 8677 2496
rect 7524 2456 7530 2468
rect 8665 2465 8677 2468
rect 8711 2465 8723 2499
rect 8665 2459 8723 2465
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7340 2400 7389 2428
rect 7340 2388 7346 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7377 2391 7435 2397
rect 7484 2400 8217 2428
rect 5997 2363 6055 2369
rect 5997 2360 6009 2363
rect 5368 2332 6009 2360
rect 5828 2304 5856 2332
rect 5997 2329 6009 2332
rect 6043 2329 6055 2363
rect 5997 2323 6055 2329
rect 6181 2363 6239 2369
rect 6181 2329 6193 2363
rect 6227 2360 6239 2363
rect 6822 2360 6828 2372
rect 6227 2332 6828 2360
rect 6227 2329 6239 2332
rect 6181 2323 6239 2329
rect 6822 2320 6828 2332
rect 6880 2360 6886 2372
rect 7484 2360 7512 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 6880 2332 7512 2360
rect 8113 2363 8171 2369
rect 6880 2320 6886 2332
rect 8113 2329 8125 2363
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 4062 2292 4068 2304
rect 3007 2264 4068 2292
rect 3007 2261 3019 2264
rect 2961 2255 3019 2261
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 5810 2252 5816 2304
rect 5868 2252 5874 2304
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 8128 2292 8156 2323
rect 6328 2264 8156 2292
rect 6328 2252 6334 2264
rect 1104 2202 9016 2224
rect 1104 2150 2599 2202
rect 2651 2150 2663 2202
rect 2715 2150 2727 2202
rect 2779 2150 2791 2202
rect 2843 2150 2855 2202
rect 2907 2150 4577 2202
rect 4629 2150 4641 2202
rect 4693 2150 4705 2202
rect 4757 2150 4769 2202
rect 4821 2150 4833 2202
rect 4885 2150 6555 2202
rect 6607 2150 6619 2202
rect 6671 2150 6683 2202
rect 6735 2150 6747 2202
rect 6799 2150 6811 2202
rect 6863 2150 8533 2202
rect 8585 2150 8597 2202
rect 8649 2150 8661 2202
rect 8713 2150 8725 2202
rect 8777 2150 8789 2202
rect 8841 2150 9016 2202
rect 1104 2128 9016 2150
rect 2958 1980 2964 2032
rect 3016 2020 3022 2032
rect 5994 2020 6000 2032
rect 3016 1992 6000 2020
rect 3016 1980 3022 1992
rect 5994 1980 6000 1992
rect 6052 1980 6058 2032
rect 1854 1912 1860 1964
rect 1912 1952 1918 1964
rect 5534 1952 5540 1964
rect 1912 1924 5540 1952
rect 1912 1912 1918 1924
rect 5534 1912 5540 1924
rect 5592 1912 5598 1964
<< via1 >>
rect 2599 9766 2651 9818
rect 2663 9766 2715 9818
rect 2727 9766 2779 9818
rect 2791 9766 2843 9818
rect 2855 9766 2907 9818
rect 4577 9766 4629 9818
rect 4641 9766 4693 9818
rect 4705 9766 4757 9818
rect 4769 9766 4821 9818
rect 4833 9766 4885 9818
rect 6555 9766 6607 9818
rect 6619 9766 6671 9818
rect 6683 9766 6735 9818
rect 6747 9766 6799 9818
rect 6811 9766 6863 9818
rect 8533 9766 8585 9818
rect 8597 9766 8649 9818
rect 8661 9766 8713 9818
rect 8725 9766 8777 9818
rect 8789 9766 8841 9818
rect 1032 9596 1084 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2964 9596 3016 9648
rect 4436 9596 4488 9648
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3792 9528 3844 9580
rect 5172 9596 5224 9648
rect 5816 9596 5868 9648
rect 4988 9528 5040 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7564 9528 7616 9580
rect 2412 9460 2464 9512
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 6644 9460 6696 9512
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8944 9528 8996 9580
rect 4344 9392 4396 9444
rect 8392 9392 8444 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 1676 9324 1728 9376
rect 2596 9324 2648 9376
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 3608 9324 3660 9376
rect 5632 9324 5684 9376
rect 6736 9324 6788 9376
rect 7380 9324 7432 9376
rect 8300 9324 8352 9376
rect 1939 9222 1991 9274
rect 2003 9222 2055 9274
rect 2067 9222 2119 9274
rect 2131 9222 2183 9274
rect 2195 9222 2247 9274
rect 3917 9222 3969 9274
rect 3981 9222 4033 9274
rect 4045 9222 4097 9274
rect 4109 9222 4161 9274
rect 4173 9222 4225 9274
rect 5895 9222 5947 9274
rect 5959 9222 6011 9274
rect 6023 9222 6075 9274
rect 6087 9222 6139 9274
rect 6151 9222 6203 9274
rect 7873 9222 7925 9274
rect 7937 9222 7989 9274
rect 8001 9222 8053 9274
rect 8065 9222 8117 9274
rect 8129 9222 8181 9274
rect 1860 9052 1912 9104
rect 3240 9120 3292 9172
rect 4344 9120 4396 9172
rect 3516 9052 3568 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 1952 8984 2004 9036
rect 3056 8984 3108 9036
rect 3608 9027 3660 9036
rect 3608 8993 3617 9027
rect 3617 8993 3651 9027
rect 3651 8993 3660 9027
rect 3608 8984 3660 8993
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2228 8848 2280 8900
rect 2596 8891 2648 8900
rect 2596 8857 2605 8891
rect 2605 8857 2639 8891
rect 2639 8857 2648 8891
rect 3424 8916 3476 8968
rect 2596 8848 2648 8857
rect 3332 8848 3384 8900
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 3700 8848 3752 8900
rect 4436 8916 4488 8968
rect 5172 9052 5224 9104
rect 7564 9120 7616 9172
rect 6368 9052 6420 9104
rect 5264 8984 5316 9036
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 8024 8984 8076 9036
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 6736 8916 6788 8968
rect 1768 8780 1820 8832
rect 1860 8780 1912 8832
rect 3056 8780 3108 8832
rect 3424 8780 3476 8832
rect 5080 8848 5132 8900
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 4252 8780 4304 8832
rect 6000 8780 6052 8832
rect 6184 8780 6236 8832
rect 8392 8959 8444 8968
rect 8392 8925 8427 8959
rect 8427 8925 8444 8959
rect 8392 8916 8444 8925
rect 8208 8891 8260 8900
rect 8208 8857 8217 8891
rect 8217 8857 8251 8891
rect 8251 8857 8260 8891
rect 8208 8848 8260 8857
rect 9036 8848 9088 8900
rect 8392 8780 8444 8832
rect 2599 8678 2651 8730
rect 2663 8678 2715 8730
rect 2727 8678 2779 8730
rect 2791 8678 2843 8730
rect 2855 8678 2907 8730
rect 4577 8678 4629 8730
rect 4641 8678 4693 8730
rect 4705 8678 4757 8730
rect 4769 8678 4821 8730
rect 4833 8678 4885 8730
rect 6555 8678 6607 8730
rect 6619 8678 6671 8730
rect 6683 8678 6735 8730
rect 6747 8678 6799 8730
rect 6811 8678 6863 8730
rect 8533 8678 8585 8730
rect 8597 8678 8649 8730
rect 8661 8678 8713 8730
rect 8725 8678 8777 8730
rect 8789 8678 8841 8730
rect 2504 8576 2556 8628
rect 2872 8619 2924 8628
rect 2872 8585 2897 8619
rect 2897 8585 2924 8619
rect 2872 8576 2924 8585
rect 3148 8576 3200 8628
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2688 8551 2740 8560
rect 2688 8517 2697 8551
rect 2697 8517 2731 8551
rect 2731 8517 2740 8551
rect 2688 8508 2740 8517
rect 3240 8551 3292 8560
rect 3240 8517 3249 8551
rect 3249 8517 3283 8551
rect 3283 8517 3292 8551
rect 3240 8508 3292 8517
rect 3700 8508 3752 8560
rect 4988 8576 5040 8628
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5448 8576 5500 8628
rect 7656 8576 7708 8628
rect 3056 8440 3108 8492
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 2688 8372 2740 8424
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 3516 8440 3568 8492
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 5080 8440 5132 8492
rect 5540 8508 5592 8560
rect 5632 8551 5684 8560
rect 5632 8517 5641 8551
rect 5641 8517 5675 8551
rect 5675 8517 5684 8551
rect 5632 8508 5684 8517
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 8300 8508 8352 8560
rect 7564 8440 7616 8492
rect 7748 8440 7800 8492
rect 8024 8372 8076 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 2320 8304 2372 8356
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 2964 8304 3016 8356
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 4896 8304 4948 8356
rect 8300 8415 8352 8424
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 9036 8372 9088 8424
rect 9128 8304 9180 8356
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 7656 8236 7708 8288
rect 8116 8236 8168 8288
rect 1939 8134 1991 8186
rect 2003 8134 2055 8186
rect 2067 8134 2119 8186
rect 2131 8134 2183 8186
rect 2195 8134 2247 8186
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 5895 8134 5947 8186
rect 5959 8134 6011 8186
rect 6023 8134 6075 8186
rect 6087 8134 6139 8186
rect 6151 8134 6203 8186
rect 7873 8134 7925 8186
rect 7937 8134 7989 8186
rect 8001 8134 8053 8186
rect 8065 8134 8117 8186
rect 8129 8134 8181 8186
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 7748 8032 7800 8084
rect 1308 7896 1360 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 3056 7896 3108 7948
rect 4436 7896 4488 7948
rect 4252 7828 4304 7880
rect 5816 7896 5868 7948
rect 6276 7896 6328 7948
rect 6920 7896 6972 7948
rect 7380 7896 7432 7948
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 7748 7939 7800 7948
rect 7748 7905 7758 7939
rect 7758 7905 7792 7939
rect 7792 7905 7800 7939
rect 7748 7896 7800 7905
rect 1400 7760 1452 7812
rect 2504 7760 2556 7812
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5356 7828 5408 7880
rect 4988 7803 5040 7812
rect 4988 7769 4997 7803
rect 4997 7769 5031 7803
rect 5031 7769 5040 7803
rect 4988 7760 5040 7769
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 1676 7692 1728 7744
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 4252 7692 4304 7744
rect 5448 7760 5500 7812
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 6276 7760 6328 7812
rect 7840 7828 7892 7880
rect 8208 7828 8260 7880
rect 8300 7828 8352 7880
rect 7012 7692 7064 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 7656 7692 7708 7744
rect 8208 7692 8260 7744
rect 8944 7692 8996 7744
rect 2599 7590 2651 7642
rect 2663 7590 2715 7642
rect 2727 7590 2779 7642
rect 2791 7590 2843 7642
rect 2855 7590 2907 7642
rect 4577 7590 4629 7642
rect 4641 7590 4693 7642
rect 4705 7590 4757 7642
rect 4769 7590 4821 7642
rect 4833 7590 4885 7642
rect 6555 7590 6607 7642
rect 6619 7590 6671 7642
rect 6683 7590 6735 7642
rect 6747 7590 6799 7642
rect 6811 7590 6863 7642
rect 8533 7590 8585 7642
rect 8597 7590 8649 7642
rect 8661 7590 8713 7642
rect 8725 7590 8777 7642
rect 8789 7590 8841 7642
rect 1860 7488 1912 7540
rect 2412 7488 2464 7540
rect 5264 7488 5316 7540
rect 5448 7488 5500 7540
rect 1676 7420 1728 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 1492 7284 1544 7336
rect 1768 7284 1820 7336
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 7196 7488 7248 7540
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 6920 7352 6972 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7840 7420 7892 7472
rect 4528 7284 4580 7336
rect 4988 7284 5040 7336
rect 8300 7352 8352 7404
rect 8484 7352 8536 7404
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 7564 7284 7616 7336
rect 7472 7216 7524 7268
rect 8392 7148 8444 7200
rect 1939 7046 1991 7098
rect 2003 7046 2055 7098
rect 2067 7046 2119 7098
rect 2131 7046 2183 7098
rect 2195 7046 2247 7098
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 5895 7046 5947 7098
rect 5959 7046 6011 7098
rect 6023 7046 6075 7098
rect 6087 7046 6139 7098
rect 6151 7046 6203 7098
rect 7873 7046 7925 7098
rect 7937 7046 7989 7098
rect 8001 7046 8053 7098
rect 8065 7046 8117 7098
rect 8129 7046 8181 7098
rect 4160 6944 4212 6996
rect 4344 6944 4396 6996
rect 5908 6944 5960 6996
rect 7104 6944 7156 6996
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 848 6604 900 6656
rect 2228 6740 2280 6792
rect 2320 6715 2372 6724
rect 2320 6681 2329 6715
rect 2329 6681 2363 6715
rect 2363 6681 2372 6715
rect 2320 6672 2372 6681
rect 2412 6672 2464 6724
rect 2964 6672 3016 6724
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 1860 6604 1912 6656
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4068 6672 4120 6724
rect 5448 6876 5500 6928
rect 6460 6876 6512 6928
rect 6920 6876 6972 6928
rect 6368 6740 6420 6792
rect 5080 6672 5132 6724
rect 5356 6672 5408 6724
rect 5816 6672 5868 6724
rect 7196 6740 7248 6792
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 7472 6740 7524 6792
rect 8116 6740 8168 6792
rect 4252 6604 4304 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 4620 6604 4672 6656
rect 5724 6604 5776 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 6000 6604 6052 6656
rect 7104 6672 7156 6724
rect 7564 6672 7616 6724
rect 8944 6672 8996 6724
rect 9128 6672 9180 6724
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 7012 6604 7064 6656
rect 8484 6604 8536 6656
rect 2599 6502 2651 6554
rect 2663 6502 2715 6554
rect 2727 6502 2779 6554
rect 2791 6502 2843 6554
rect 2855 6502 2907 6554
rect 4577 6502 4629 6554
rect 4641 6502 4693 6554
rect 4705 6502 4757 6554
rect 4769 6502 4821 6554
rect 4833 6502 4885 6554
rect 6555 6502 6607 6554
rect 6619 6502 6671 6554
rect 6683 6502 6735 6554
rect 6747 6502 6799 6554
rect 6811 6502 6863 6554
rect 8533 6502 8585 6554
rect 8597 6502 8649 6554
rect 8661 6502 8713 6554
rect 8725 6502 8777 6554
rect 8789 6502 8841 6554
rect 2320 6400 2372 6452
rect 2596 6400 2648 6452
rect 1400 6332 1452 6384
rect 4068 6400 4120 6452
rect 6276 6400 6328 6452
rect 6644 6400 6696 6452
rect 8116 6400 8168 6452
rect 8484 6400 8536 6452
rect 9036 6400 9088 6452
rect 2136 6264 2188 6316
rect 2504 6264 2556 6316
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 3148 6332 3200 6384
rect 2780 6264 2832 6273
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 4344 6264 4396 6316
rect 4988 6332 5040 6384
rect 7104 6332 7156 6384
rect 2504 6128 2556 6180
rect 1676 6060 1728 6112
rect 1768 6060 1820 6112
rect 3056 6128 3108 6180
rect 4252 6196 4304 6248
rect 5356 6264 5408 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6920 6264 6972 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 2780 6060 2832 6112
rect 3516 6060 3568 6112
rect 5632 6196 5684 6248
rect 6276 6196 6328 6248
rect 4896 6060 4948 6112
rect 4988 6060 5040 6112
rect 6368 6128 6420 6180
rect 7012 6060 7064 6112
rect 7656 6060 7708 6112
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 1939 5958 1991 6010
rect 2003 5958 2055 6010
rect 2067 5958 2119 6010
rect 2131 5958 2183 6010
rect 2195 5958 2247 6010
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 5895 5958 5947 6010
rect 5959 5958 6011 6010
rect 6023 5958 6075 6010
rect 6087 5958 6139 6010
rect 6151 5958 6203 6010
rect 7873 5958 7925 6010
rect 7937 5958 7989 6010
rect 8001 5958 8053 6010
rect 8065 5958 8117 6010
rect 8129 5958 8181 6010
rect 3516 5856 3568 5908
rect 3608 5856 3660 5908
rect 4252 5856 4304 5908
rect 5172 5856 5224 5908
rect 5724 5856 5776 5908
rect 5908 5856 5960 5908
rect 7380 5856 7432 5908
rect 2412 5788 2464 5840
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 1860 5720 1912 5772
rect 848 5652 900 5704
rect 1492 5652 1544 5704
rect 5816 5788 5868 5840
rect 7932 5788 7984 5840
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 7472 5720 7524 5772
rect 7748 5720 7800 5772
rect 8944 5788 8996 5840
rect 1768 5584 1820 5636
rect 1952 5627 2004 5636
rect 1952 5593 1961 5627
rect 1961 5593 1995 5627
rect 1995 5593 2004 5627
rect 1952 5584 2004 5593
rect 3148 5584 3200 5636
rect 2412 5516 2464 5568
rect 2688 5516 2740 5568
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 4252 5584 4304 5636
rect 5356 5652 5408 5704
rect 6368 5652 6420 5704
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 4896 5584 4948 5636
rect 5448 5627 5500 5636
rect 5448 5593 5457 5627
rect 5457 5593 5491 5627
rect 5491 5593 5500 5627
rect 5448 5584 5500 5593
rect 5540 5584 5592 5636
rect 5908 5627 5960 5636
rect 5908 5593 5917 5627
rect 5917 5593 5951 5627
rect 5951 5593 5960 5627
rect 5908 5584 5960 5593
rect 7104 5652 7156 5704
rect 7380 5652 7432 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 6920 5627 6972 5636
rect 6920 5593 6929 5627
rect 6929 5593 6963 5627
rect 6963 5593 6972 5627
rect 6920 5584 6972 5593
rect 7472 5584 7524 5636
rect 8392 5584 8444 5636
rect 3424 5516 3476 5568
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 6000 5516 6052 5568
rect 6184 5516 6236 5568
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 8208 5516 8260 5568
rect 8484 5516 8536 5568
rect 2599 5414 2651 5466
rect 2663 5414 2715 5466
rect 2727 5414 2779 5466
rect 2791 5414 2843 5466
rect 2855 5414 2907 5466
rect 4577 5414 4629 5466
rect 4641 5414 4693 5466
rect 4705 5414 4757 5466
rect 4769 5414 4821 5466
rect 4833 5414 4885 5466
rect 6555 5414 6607 5466
rect 6619 5414 6671 5466
rect 6683 5414 6735 5466
rect 6747 5414 6799 5466
rect 6811 5414 6863 5466
rect 8533 5414 8585 5466
rect 8597 5414 8649 5466
rect 8661 5414 8713 5466
rect 8725 5414 8777 5466
rect 8789 5414 8841 5466
rect 2412 5312 2464 5364
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 5632 5312 5684 5364
rect 940 5244 992 5296
rect 2320 5176 2372 5228
rect 3792 5244 3844 5296
rect 4804 5287 4856 5296
rect 4804 5253 4813 5287
rect 4813 5253 4847 5287
rect 4847 5253 4856 5287
rect 4804 5244 4856 5253
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 4344 5176 4396 5228
rect 4620 5176 4672 5228
rect 2504 5108 2556 5160
rect 5080 5176 5132 5228
rect 4988 5108 5040 5160
rect 5632 5219 5684 5229
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5177 5684 5185
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 6092 5312 6144 5364
rect 6000 5244 6052 5296
rect 6184 5176 6236 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6736 5176 6788 5228
rect 6828 5108 6880 5160
rect 5448 5040 5500 5092
rect 6920 5040 6972 5092
rect 7288 5040 7340 5092
rect 7380 5083 7432 5092
rect 7380 5049 7389 5083
rect 7389 5049 7423 5083
rect 7423 5049 7432 5083
rect 7380 5040 7432 5049
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 3148 4972 3200 4981
rect 3700 4972 3752 5024
rect 8392 4972 8444 5024
rect 1939 4870 1991 4922
rect 2003 4870 2055 4922
rect 2067 4870 2119 4922
rect 2131 4870 2183 4922
rect 2195 4870 2247 4922
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 5895 4870 5947 4922
rect 5959 4870 6011 4922
rect 6023 4870 6075 4922
rect 6087 4870 6139 4922
rect 6151 4870 6203 4922
rect 7873 4870 7925 4922
rect 7937 4870 7989 4922
rect 8001 4870 8053 4922
rect 8065 4870 8117 4922
rect 8129 4870 8181 4922
rect 4160 4768 4212 4820
rect 4620 4768 4672 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 8300 4768 8352 4820
rect 2504 4632 2556 4684
rect 2964 4700 3016 4752
rect 4804 4700 4856 4752
rect 5264 4743 5316 4752
rect 5264 4709 5273 4743
rect 5273 4709 5307 4743
rect 5307 4709 5316 4743
rect 5264 4700 5316 4709
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 5172 4632 5224 4684
rect 5816 4632 5868 4684
rect 1400 4564 1452 4616
rect 2964 4564 3016 4616
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 7196 4632 7248 4684
rect 7656 4632 7708 4684
rect 7748 4564 7800 4616
rect 2412 4496 2464 4548
rect 3608 4496 3660 4548
rect 4896 4496 4948 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2044 4471 2096 4480
rect 2044 4437 2053 4471
rect 2053 4437 2087 4471
rect 2087 4437 2096 4471
rect 2044 4428 2096 4437
rect 3792 4428 3844 4480
rect 5080 4496 5132 4548
rect 5724 4428 5776 4480
rect 2599 4326 2651 4378
rect 2663 4326 2715 4378
rect 2727 4326 2779 4378
rect 2791 4326 2843 4378
rect 2855 4326 2907 4378
rect 4577 4326 4629 4378
rect 4641 4326 4693 4378
rect 4705 4326 4757 4378
rect 4769 4326 4821 4378
rect 4833 4326 4885 4378
rect 6555 4326 6607 4378
rect 6619 4326 6671 4378
rect 6683 4326 6735 4378
rect 6747 4326 6799 4378
rect 6811 4326 6863 4378
rect 8533 4326 8585 4378
rect 8597 4326 8649 4378
rect 8661 4326 8713 4378
rect 8725 4326 8777 4378
rect 8789 4326 8841 4378
rect 2044 4224 2096 4276
rect 2320 4224 2372 4276
rect 2412 4224 2464 4276
rect 3240 4224 3292 4276
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 1768 3952 1820 4004
rect 2504 4088 2556 4140
rect 2780 4156 2832 4208
rect 3608 4156 3660 4208
rect 4252 4267 4304 4276
rect 4252 4233 4261 4267
rect 4261 4233 4295 4267
rect 4295 4233 4304 4267
rect 4252 4224 4304 4233
rect 4436 4224 4488 4276
rect 5632 4224 5684 4276
rect 7104 4224 7156 4276
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 3056 4088 3108 4140
rect 3608 4020 3660 4072
rect 4436 4088 4488 4140
rect 4344 4020 4396 4072
rect 5172 4156 5224 4208
rect 7196 4156 7248 4208
rect 5356 4088 5408 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 5816 4088 5868 4140
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 6368 4088 6420 4140
rect 6276 4020 6328 4072
rect 6368 3952 6420 4004
rect 6920 4020 6972 4072
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 7380 4088 7432 4140
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 7656 4063 7708 4072
rect 7656 4029 7665 4063
rect 7665 4029 7699 4063
rect 7699 4029 7708 4063
rect 7656 4020 7708 4029
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 8944 3952 8996 4004
rect 2320 3884 2372 3936
rect 3148 3884 3200 3936
rect 3332 3884 3384 3936
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 5540 3884 5592 3936
rect 1939 3782 1991 3834
rect 2003 3782 2055 3834
rect 2067 3782 2119 3834
rect 2131 3782 2183 3834
rect 2195 3782 2247 3834
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 5895 3782 5947 3834
rect 5959 3782 6011 3834
rect 6023 3782 6075 3834
rect 6087 3782 6139 3834
rect 6151 3782 6203 3834
rect 7873 3782 7925 3834
rect 7937 3782 7989 3834
rect 8001 3782 8053 3834
rect 8065 3782 8117 3834
rect 8129 3782 8181 3834
rect 1768 3680 1820 3732
rect 2412 3680 2464 3732
rect 2964 3680 3016 3732
rect 3976 3680 4028 3732
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 5632 3680 5684 3732
rect 8484 3680 8536 3732
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 3516 3544 3568 3596
rect 4068 3544 4120 3596
rect 3240 3476 3292 3528
rect 3792 3476 3844 3528
rect 4988 3544 5040 3596
rect 5264 3544 5316 3596
rect 5356 3544 5408 3596
rect 6920 3612 6972 3664
rect 7288 3612 7340 3664
rect 8208 3612 8260 3664
rect 3884 3408 3936 3460
rect 4160 3451 4212 3460
rect 4160 3417 4185 3451
rect 4185 3417 4212 3451
rect 4160 3408 4212 3417
rect 2504 3340 2556 3392
rect 2780 3340 2832 3392
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 3056 3340 3108 3392
rect 3608 3340 3660 3392
rect 4344 3340 4396 3392
rect 4528 3408 4580 3460
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 7748 3544 7800 3596
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7196 3519 7248 3528
rect 7196 3485 7205 3519
rect 7205 3485 7239 3519
rect 7239 3485 7248 3519
rect 7196 3476 7248 3485
rect 5080 3340 5132 3392
rect 5540 3340 5592 3392
rect 6368 3408 6420 3460
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 7748 3408 7800 3460
rect 8392 3408 8444 3460
rect 6828 3383 6880 3392
rect 6828 3349 6837 3383
rect 6837 3349 6871 3383
rect 6871 3349 6880 3383
rect 6828 3340 6880 3349
rect 8116 3340 8168 3392
rect 2599 3238 2651 3290
rect 2663 3238 2715 3290
rect 2727 3238 2779 3290
rect 2791 3238 2843 3290
rect 2855 3238 2907 3290
rect 4577 3238 4629 3290
rect 4641 3238 4693 3290
rect 4705 3238 4757 3290
rect 4769 3238 4821 3290
rect 4833 3238 4885 3290
rect 6555 3238 6607 3290
rect 6619 3238 6671 3290
rect 6683 3238 6735 3290
rect 6747 3238 6799 3290
rect 6811 3238 6863 3290
rect 8533 3238 8585 3290
rect 8597 3238 8649 3290
rect 8661 3238 8713 3290
rect 8725 3238 8777 3290
rect 8789 3238 8841 3290
rect 1860 3136 1912 3188
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 2412 3068 2464 3120
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 1768 3000 1820 3052
rect 1860 3000 1912 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 1952 2932 2004 2984
rect 2964 3068 3016 3120
rect 3424 3136 3476 3188
rect 3608 3136 3660 3188
rect 3884 3068 3936 3120
rect 4068 3068 4120 3120
rect 4436 3136 4488 3188
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 6644 3136 6696 3188
rect 7380 3136 7432 3188
rect 7472 3136 7524 3188
rect 7840 3136 7892 3188
rect 8300 3136 8352 3188
rect 5172 3068 5224 3120
rect 4344 3000 4396 3052
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5632 3000 5684 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8208 3000 8260 3052
rect 6828 2932 6880 2984
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 2596 2864 2648 2916
rect 4160 2864 4212 2916
rect 4436 2864 4488 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 2320 2796 2372 2848
rect 3516 2796 3568 2848
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 5724 2839 5776 2848
rect 5724 2805 5733 2839
rect 5733 2805 5767 2839
rect 5767 2805 5776 2839
rect 5724 2796 5776 2805
rect 6460 2796 6512 2848
rect 7196 2796 7248 2848
rect 7288 2796 7340 2848
rect 7840 2932 7892 2984
rect 7748 2864 7800 2916
rect 8300 2796 8352 2848
rect 1939 2694 1991 2746
rect 2003 2694 2055 2746
rect 2067 2694 2119 2746
rect 2131 2694 2183 2746
rect 2195 2694 2247 2746
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 5895 2694 5947 2746
rect 5959 2694 6011 2746
rect 6023 2694 6075 2746
rect 6087 2694 6139 2746
rect 6151 2694 6203 2746
rect 7873 2694 7925 2746
rect 7937 2694 7989 2746
rect 8001 2694 8053 2746
rect 8065 2694 8117 2746
rect 8129 2694 8181 2746
rect 1584 2592 1636 2644
rect 2228 2592 2280 2644
rect 2412 2592 2464 2644
rect 2412 2456 2464 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 3056 2592 3108 2644
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4436 2592 4488 2644
rect 5540 2592 5592 2644
rect 6276 2592 6328 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 2596 2567 2648 2576
rect 2596 2533 2605 2567
rect 2605 2533 2639 2567
rect 2639 2533 2648 2567
rect 2596 2524 2648 2533
rect 5264 2524 5316 2576
rect 5448 2524 5500 2576
rect 7012 2592 7064 2644
rect 7380 2592 7432 2644
rect 7564 2592 7616 2644
rect 8392 2592 8444 2644
rect 2872 2388 2924 2440
rect 1768 2320 1820 2372
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 1860 2252 1912 2261
rect 2320 2252 2372 2304
rect 5540 2456 5592 2508
rect 3424 2388 3476 2440
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 3700 2388 3752 2440
rect 4160 2388 4212 2440
rect 4436 2363 4488 2372
rect 4436 2329 4445 2363
rect 4445 2329 4479 2363
rect 4479 2329 4488 2363
rect 4436 2320 4488 2329
rect 5172 2320 5224 2372
rect 5724 2388 5776 2440
rect 7472 2456 7524 2508
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7288 2388 7340 2440
rect 6828 2320 6880 2372
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 4068 2252 4120 2304
rect 5816 2252 5868 2304
rect 6276 2252 6328 2304
rect 2599 2150 2651 2202
rect 2663 2150 2715 2202
rect 2727 2150 2779 2202
rect 2791 2150 2843 2202
rect 2855 2150 2907 2202
rect 4577 2150 4629 2202
rect 4641 2150 4693 2202
rect 4705 2150 4757 2202
rect 4769 2150 4821 2202
rect 4833 2150 4885 2202
rect 6555 2150 6607 2202
rect 6619 2150 6671 2202
rect 6683 2150 6735 2202
rect 6747 2150 6799 2202
rect 6811 2150 6863 2202
rect 8533 2150 8585 2202
rect 8597 2150 8649 2202
rect 8661 2150 8713 2202
rect 8725 2150 8777 2202
rect 8789 2150 8841 2202
rect 2964 1980 3016 2032
rect 6000 1980 6052 2032
rect 1860 1912 1912 1964
rect 5540 1912 5592 1964
<< metal2 >>
rect 4526 11545 4582 12345
rect 5170 11545 5226 12345
rect 5814 11545 5870 12345
rect 4540 10554 4568 11545
rect 4448 10526 4568 10554
rect 2599 9820 2907 9829
rect 2599 9818 2605 9820
rect 2661 9818 2685 9820
rect 2741 9818 2765 9820
rect 2821 9818 2845 9820
rect 2901 9818 2907 9820
rect 2661 9766 2663 9818
rect 2843 9766 2845 9818
rect 2599 9764 2605 9766
rect 2661 9764 2685 9766
rect 2741 9764 2765 9766
rect 2821 9764 2845 9766
rect 2901 9764 2907 9766
rect 2599 9755 2907 9764
rect 4448 9654 4476 10526
rect 4577 9820 4885 9829
rect 4577 9818 4583 9820
rect 4639 9818 4663 9820
rect 4719 9818 4743 9820
rect 4799 9818 4823 9820
rect 4879 9818 4885 9820
rect 4639 9766 4641 9818
rect 4821 9766 4823 9818
rect 4577 9764 4583 9766
rect 4639 9764 4663 9766
rect 4719 9764 4743 9766
rect 4799 9764 4823 9766
rect 4879 9764 4885 9766
rect 4577 9755 4885 9764
rect 5184 9654 5212 11545
rect 5828 9654 5856 11545
rect 6555 9820 6863 9829
rect 6555 9818 6561 9820
rect 6617 9818 6641 9820
rect 6697 9818 6721 9820
rect 6777 9818 6801 9820
rect 6857 9818 6863 9820
rect 6617 9766 6619 9818
rect 6799 9766 6801 9818
rect 6555 9764 6561 9766
rect 6617 9764 6641 9766
rect 6697 9764 6721 9766
rect 6777 9764 6801 9766
rect 6857 9764 6863 9766
rect 6555 9755 6863 9764
rect 8533 9820 8841 9829
rect 8533 9818 8539 9820
rect 8595 9818 8619 9820
rect 8675 9818 8699 9820
rect 8755 9818 8779 9820
rect 8835 9818 8841 9820
rect 8595 9766 8597 9818
rect 8777 9766 8779 9818
rect 8533 9764 8539 9766
rect 8595 9764 8619 9766
rect 8675 9764 8699 9766
rect 8755 9764 8779 9766
rect 8835 9764 8841 9766
rect 8533 9755 8841 9764
rect 1032 9648 1084 9654
rect 1030 9616 1032 9625
rect 2964 9648 3016 9654
rect 1084 9616 1086 9625
rect 2964 9590 3016 9596
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 1030 9551 1086 9560
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 8945 1440 9522
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1596 9042 1624 9318
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1398 8936 1454 8945
rect 1398 8871 1454 8880
rect 1688 8498 1716 9318
rect 1939 9276 2247 9285
rect 1939 9274 1945 9276
rect 2001 9274 2025 9276
rect 2081 9274 2105 9276
rect 2161 9274 2185 9276
rect 2241 9274 2247 9276
rect 2001 9222 2003 9274
rect 2183 9222 2185 9274
rect 1939 9220 1945 9222
rect 2001 9220 2025 9222
rect 2081 9220 2105 9222
rect 2161 9220 2185 9222
rect 2241 9220 2247 9222
rect 1939 9211 2247 9220
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1872 8974 1900 9046
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 1320 7585 1348 7890
rect 1400 7812 1452 7818
rect 1400 7754 1452 7760
rect 1306 7576 1362 7585
rect 1306 7511 1362 7520
rect 848 6656 900 6662
rect 846 6624 848 6633
rect 900 6624 902 6633
rect 846 6559 902 6568
rect 1412 6390 1440 7754
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1596 7410 1624 7686
rect 1688 7478 1716 7686
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1780 7342 1808 8774
rect 1872 7546 1900 8774
rect 1964 8498 1992 8978
rect 2228 8900 2280 8906
rect 2228 8842 2280 8848
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2240 8294 2268 8842
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 1939 8188 2247 8197
rect 1939 8186 1945 8188
rect 2001 8186 2025 8188
rect 2081 8186 2105 8188
rect 2161 8186 2185 8188
rect 2241 8186 2247 8188
rect 2001 8134 2003 8186
rect 2183 8134 2185 8186
rect 1939 8132 1945 8134
rect 2001 8132 2025 8134
rect 2081 8132 2105 8134
rect 2161 8132 2185 8134
rect 2241 8132 2247 8134
rect 1939 8123 2247 8132
rect 2332 7886 2360 8298
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 846 5944 902 5953
rect 846 5879 902 5888
rect 860 5710 888 5879
rect 1412 5817 1440 6326
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 952 5302 980 5471
rect 940 5296 992 5302
rect 940 5238 992 5244
rect 1412 4622 1440 5743
rect 1504 5710 1532 7278
rect 2240 7188 2268 7822
rect 2424 7546 2452 9454
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8922 2636 9318
rect 2516 8906 2636 8922
rect 2516 8900 2648 8906
rect 2516 8894 2596 8900
rect 2516 8634 2544 8894
rect 2596 8842 2648 8848
rect 2599 8732 2907 8741
rect 2599 8730 2605 8732
rect 2661 8730 2685 8732
rect 2741 8730 2765 8732
rect 2821 8730 2845 8732
rect 2901 8730 2907 8732
rect 2661 8678 2663 8730
rect 2843 8678 2845 8730
rect 2599 8676 2605 8678
rect 2661 8676 2685 8678
rect 2741 8676 2765 8678
rect 2821 8676 2845 8678
rect 2901 8676 2907 8678
rect 2599 8667 2907 8676
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2872 8628 2924 8634
rect 2976 8616 3004 9590
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 3068 9042 3096 9522
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2924 8588 3004 8616
rect 2872 8570 2924 8576
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2700 8430 2728 8502
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2976 8362 3004 8588
rect 3068 8498 3096 8774
rect 3160 8634 3188 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3252 8566 3280 9114
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3160 8378 3188 8434
rect 3344 8378 3372 8842
rect 3436 8838 3464 8910
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8498 3464 8774
rect 3528 8498 3556 9046
rect 3620 9042 3648 9318
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3804 8974 3832 9522
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 3917 9276 4225 9285
rect 3917 9274 3923 9276
rect 3979 9274 4003 9276
rect 4059 9274 4083 9276
rect 4139 9274 4163 9276
rect 4219 9274 4225 9276
rect 3979 9222 3981 9274
rect 4161 9222 4163 9274
rect 3917 9220 3923 9222
rect 3979 9220 4003 9222
rect 4059 9220 4083 9222
rect 4139 9220 4163 9222
rect 4219 9220 4225 9222
rect 3917 9211 4225 9220
rect 4356 9178 4384 9386
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3712 8566 3740 8842
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 2964 8356 3016 8362
rect 3160 8350 3372 8378
rect 2964 8298 3016 8304
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3068 7954 3096 8230
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2240 7160 2360 7188
rect 1939 7100 2247 7109
rect 1939 7098 1945 7100
rect 2001 7098 2025 7100
rect 2081 7098 2105 7100
rect 2161 7098 2185 7100
rect 2241 7098 2247 7100
rect 2001 7046 2003 7098
rect 2183 7046 2185 7098
rect 1939 7044 1945 7046
rect 2001 7044 2025 7046
rect 2081 7044 2105 7046
rect 2161 7044 2185 7046
rect 2241 7044 2247 7046
rect 1939 7035 2247 7044
rect 2332 6882 2360 7160
rect 2148 6854 2360 6882
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1688 5778 1716 6054
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1780 5642 1808 6054
rect 1872 5778 1900 6598
rect 2148 6322 2176 6854
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2240 6168 2268 6734
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2332 6458 2360 6666
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2240 6140 2360 6168
rect 1939 6012 2247 6021
rect 1939 6010 1945 6012
rect 2001 6010 2025 6012
rect 2081 6010 2105 6012
rect 2161 6010 2185 6012
rect 2241 6010 2247 6012
rect 2001 5958 2003 6010
rect 2183 5958 2185 6010
rect 1939 5956 1945 5958
rect 2001 5956 2025 5958
rect 2081 5956 2105 5958
rect 2161 5956 2185 5958
rect 2241 5956 2247 5958
rect 1939 5947 2247 5956
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 2332 5710 2360 6140
rect 2424 5846 2452 6666
rect 2516 6322 2544 7754
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2599 7644 2907 7653
rect 2599 7642 2605 7644
rect 2661 7642 2685 7644
rect 2741 7642 2765 7644
rect 2821 7642 2845 7644
rect 2901 7642 2907 7644
rect 2661 7590 2663 7642
rect 2843 7590 2845 7642
rect 2599 7588 2605 7590
rect 2661 7588 2685 7590
rect 2741 7588 2765 7590
rect 2821 7588 2845 7590
rect 2901 7588 2907 7590
rect 2599 7579 2907 7588
rect 2976 6730 3004 7686
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2599 6556 2907 6565
rect 2599 6554 2605 6556
rect 2661 6554 2685 6556
rect 2741 6554 2765 6556
rect 2821 6554 2845 6556
rect 2901 6554 2907 6556
rect 2661 6502 2663 6554
rect 2843 6502 2845 6554
rect 2599 6500 2605 6502
rect 2661 6500 2685 6502
rect 2741 6500 2765 6502
rect 2821 6500 2845 6502
rect 2901 6500 2907 6502
rect 2599 6491 2907 6500
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2504 6316 2556 6322
rect 2608 6304 2636 6394
rect 2976 6322 3004 6666
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 2780 6316 2832 6322
rect 2608 6276 2780 6304
rect 2504 6258 2556 6264
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 1768 5636 1820 5642
rect 1952 5636 2004 5642
rect 1768 5578 1820 5584
rect 1872 5596 1952 5624
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4865 1532 4966
rect 1490 4856 1546 4865
rect 1490 4791 1546 4800
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4146 1624 4422
rect 1872 4146 1900 5596
rect 1952 5578 2004 5584
rect 2424 5574 2452 5646
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5370 2452 5510
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 1939 4924 2247 4933
rect 1939 4922 1945 4924
rect 2001 4922 2025 4924
rect 2081 4922 2105 4924
rect 2161 4922 2185 4924
rect 2241 4922 2247 4924
rect 2001 4870 2003 4922
rect 2183 4870 2185 4922
rect 1939 4868 1945 4870
rect 2001 4868 2025 4870
rect 2081 4868 2105 4870
rect 2161 4868 2185 4870
rect 2241 4868 2247 4870
rect 1939 4859 2247 4868
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 2056 4282 2084 4422
rect 2332 4282 2360 5170
rect 2516 5166 2544 6122
rect 2700 5574 2728 6276
rect 2780 6258 2832 6264
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2780 6112 2832 6118
rect 2832 6072 3004 6100
rect 2780 6054 2832 6060
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2599 5468 2907 5477
rect 2599 5466 2605 5468
rect 2661 5466 2685 5468
rect 2741 5466 2765 5468
rect 2821 5466 2845 5468
rect 2901 5466 2907 5468
rect 2661 5414 2663 5466
rect 2843 5414 2845 5466
rect 2599 5412 2605 5414
rect 2661 5412 2685 5414
rect 2741 5412 2765 5414
rect 2821 5412 2845 5414
rect 2901 5412 2907 5414
rect 2599 5403 2907 5412
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2516 4690 2544 5102
rect 2976 4758 3004 6072
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2424 4282 2452 4490
rect 2599 4380 2907 4389
rect 2599 4378 2605 4380
rect 2661 4378 2685 4380
rect 2741 4378 2765 4380
rect 2821 4378 2845 4380
rect 2901 4378 2907 4380
rect 2661 4326 2663 4378
rect 2843 4326 2845 4378
rect 2599 4324 2605 4326
rect 2661 4324 2685 4326
rect 2741 4324 2765 4326
rect 2821 4324 2845 4326
rect 2901 4324 2907 4326
rect 2599 4315 2907 4324
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1964 4026 1992 4082
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 1872 3998 1992 4026
rect 1780 3738 1808 3946
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1676 3528 1728 3534
rect 1452 3496 1454 3505
rect 1676 3470 1728 3476
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1398 3431 1454 3440
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1596 2650 1624 2994
rect 1688 2854 1716 3470
rect 1780 3058 1808 3470
rect 1872 3194 1900 3998
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1939 3836 2247 3845
rect 1939 3834 1945 3836
rect 2001 3834 2025 3836
rect 2081 3834 2105 3836
rect 2161 3834 2185 3836
rect 2241 3834 2247 3836
rect 2001 3782 2003 3834
rect 2183 3782 2185 3834
rect 1939 3780 1945 3782
rect 2001 3780 2025 3782
rect 2081 3780 2105 3782
rect 2161 3780 2185 3782
rect 2241 3780 2247 3782
rect 1939 3771 2247 3780
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1872 2774 1900 2994
rect 1964 2990 1992 3538
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 3126 2084 3470
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2332 2854 2360 3878
rect 2424 3738 2452 4218
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2516 3482 2544 4082
rect 2424 3454 2544 3482
rect 2424 3126 2452 3454
rect 2792 3398 2820 4150
rect 2976 3738 3004 4558
rect 3068 4146 3096 6122
rect 3160 5642 3188 6326
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5914 3556 6054
rect 3620 5914 3648 6598
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3148 5636 3200 5642
rect 3200 5596 3280 5624
rect 3148 5578 3200 5584
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3160 4026 3188 4966
rect 3252 4282 3280 5596
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 5234 3464 5510
rect 3620 5234 3648 5850
rect 3712 5234 3740 8502
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 4264 7886 4292 8774
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4172 6798 4200 6938
rect 4264 6798 4292 7686
rect 4356 7002 4384 8230
rect 4448 7954 4476 8910
rect 4577 8732 4885 8741
rect 4577 8730 4583 8732
rect 4639 8730 4663 8732
rect 4719 8730 4743 8732
rect 4799 8730 4823 8732
rect 4879 8730 4885 8732
rect 4639 8678 4641 8730
rect 4821 8678 4823 8730
rect 4577 8676 4583 8678
rect 4639 8676 4663 8678
rect 4719 8676 4743 8678
rect 4799 8676 4823 8678
rect 4879 8676 4885 8678
rect 4577 8667 4885 8676
rect 5000 8634 5028 9522
rect 5092 8906 5120 9522
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5092 8498 5120 8842
rect 5184 8634 5212 9046
rect 5276 9042 5304 9454
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4632 8090 4660 8434
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 5710 3832 6598
rect 4080 6458 4108 6666
rect 4264 6662 4292 6734
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4356 6322 4384 6598
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4252 6248 4304 6254
rect 4448 6202 4476 7890
rect 4908 7886 4936 8298
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4577 7644 4885 7653
rect 4577 7642 4583 7644
rect 4639 7642 4663 7644
rect 4719 7642 4743 7644
rect 4799 7642 4823 7644
rect 4879 7642 4885 7644
rect 4639 7590 4641 7642
rect 4821 7590 4823 7642
rect 4577 7588 4583 7590
rect 4639 7588 4663 7590
rect 4719 7588 4743 7590
rect 4799 7588 4823 7590
rect 4879 7588 4885 7590
rect 4577 7579 4885 7588
rect 5000 7342 5028 7754
rect 5276 7546 5304 7822
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4988 7336 5040 7342
rect 5368 7313 5396 7822
rect 5460 7818 5488 8570
rect 5552 8566 5580 8910
rect 5644 8566 5672 9318
rect 5895 9276 6203 9285
rect 5895 9274 5901 9276
rect 5957 9274 5981 9276
rect 6037 9274 6061 9276
rect 6117 9274 6141 9276
rect 6197 9274 6203 9276
rect 5957 9222 5959 9274
rect 6139 9222 6141 9274
rect 5895 9220 5901 9222
rect 5957 9220 5981 9222
rect 6037 9220 6061 9222
rect 6117 9220 6141 9222
rect 6197 9220 6203 9222
rect 5895 9211 6203 9220
rect 6380 9110 6408 9454
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6656 9042 6684 9454
rect 6748 9382 6776 9522
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6748 8974 6776 9318
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7010 8936 7066 8945
rect 7010 8871 7066 8880
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5632 8560 5684 8566
rect 5632 8502 5684 8508
rect 6012 8498 6040 8774
rect 6196 8498 6224 8774
rect 6555 8732 6863 8741
rect 6555 8730 6561 8732
rect 6617 8730 6641 8732
rect 6697 8730 6721 8732
rect 6777 8730 6801 8732
rect 6857 8730 6863 8732
rect 6617 8678 6619 8730
rect 6799 8678 6801 8730
rect 6555 8676 6561 8678
rect 6617 8676 6641 8678
rect 6697 8676 6721 8678
rect 6777 8676 6801 8678
rect 6857 8676 6863 8678
rect 6555 8667 6863 8676
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6196 8344 6224 8434
rect 6196 8316 6316 8344
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5828 7954 5856 8230
rect 5895 8188 6203 8197
rect 5895 8186 5901 8188
rect 5957 8186 5981 8188
rect 6037 8186 6061 8188
rect 6117 8186 6141 8188
rect 6197 8186 6203 8188
rect 5957 8134 5959 8186
rect 6139 8134 6141 8186
rect 5895 8132 5901 8134
rect 5957 8132 5981 8134
rect 6037 8132 6061 8134
rect 6117 8132 6141 8134
rect 6197 8132 6203 8134
rect 5895 8123 6203 8132
rect 6288 7954 6316 8316
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 5460 7546 5488 7754
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 4988 7278 5040 7284
rect 5354 7304 5410 7313
rect 4540 6644 4568 7278
rect 4620 6656 4672 6662
rect 4508 6616 4620 6644
rect 4508 6440 4536 6616
rect 4620 6598 4672 6604
rect 4577 6556 4885 6565
rect 4577 6554 4583 6556
rect 4639 6554 4663 6556
rect 4719 6554 4743 6556
rect 4799 6554 4823 6556
rect 4879 6554 4885 6556
rect 4639 6502 4641 6554
rect 4821 6502 4823 6554
rect 4577 6500 4583 6502
rect 4639 6500 4663 6502
rect 4719 6500 4743 6502
rect 4799 6500 4823 6502
rect 4879 6500 4885 6502
rect 4577 6491 4885 6500
rect 4508 6412 4568 6440
rect 4304 6196 4476 6202
rect 4252 6190 4476 6196
rect 4264 6174 4476 6190
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 4264 5914 4292 6174
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4342 5808 4398 5817
rect 4540 5794 4568 6412
rect 5000 6390 5028 7278
rect 5354 7239 5410 7248
rect 5368 6730 5396 7239
rect 5460 6934 5488 7346
rect 5895 7100 6203 7109
rect 5895 7098 5901 7100
rect 5957 7098 5981 7100
rect 6037 7098 6061 7100
rect 6117 7098 6141 7100
rect 6197 7098 6203 7100
rect 5957 7046 5959 7098
rect 6139 7046 6141 7098
rect 5895 7044 5901 7046
rect 5957 7044 5981 7046
rect 6037 7044 6061 7046
rect 6117 7044 6141 7046
rect 6197 7044 6203 7046
rect 5895 7035 6203 7044
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 4988 6384 5040 6390
rect 4988 6326 5040 6332
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4398 5766 4568 5794
rect 4342 5743 4344 5752
rect 4396 5743 4398 5752
rect 4344 5714 4396 5720
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 3804 5302 3832 5646
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5370 4292 5578
rect 4252 5364 4304 5370
rect 4448 5352 4476 5646
rect 4908 5642 4936 6054
rect 4896 5636 4948 5642
rect 4896 5578 4948 5584
rect 4577 5468 4885 5477
rect 4577 5466 4583 5468
rect 4639 5466 4663 5468
rect 4719 5466 4743 5468
rect 4799 5466 4823 5468
rect 4879 5466 4885 5468
rect 4639 5414 4641 5466
rect 4821 5414 4823 5466
rect 4577 5412 4583 5414
rect 4639 5412 4663 5414
rect 4719 5412 4743 5414
rect 4799 5412 4823 5414
rect 4879 5412 4885 5414
rect 4577 5403 4885 5412
rect 5000 5386 5028 6054
rect 5092 5681 5120 6666
rect 5368 6322 5396 6666
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6322 5764 6598
rect 5828 6322 5856 6666
rect 5920 6662 5948 6938
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5078 5672 5134 5681
rect 5078 5607 5134 5616
rect 5092 5574 5120 5607
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4908 5358 5028 5386
rect 4448 5324 4660 5352
rect 4252 5306 4304 5312
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 4632 5234 4660 5324
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 4344 5228 4396 5234
rect 4620 5228 4672 5234
rect 4396 5188 4476 5216
rect 4344 5170 4396 5176
rect 3712 5114 3740 5170
rect 3620 5086 3740 5114
rect 3620 4554 3648 5086
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3620 4214 3648 4490
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3608 4072 3660 4078
rect 3160 3998 3464 4026
rect 3608 4014 3660 4020
rect 3160 3942 3188 3998
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1780 2746 1900 2774
rect 1939 2748 2247 2757
rect 1939 2746 1945 2748
rect 2001 2746 2025 2748
rect 2081 2746 2105 2748
rect 2161 2746 2185 2748
rect 2241 2746 2247 2748
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 1688 2446 1716 2479
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1780 2378 1808 2746
rect 2001 2694 2003 2746
rect 2183 2694 2185 2746
rect 1939 2692 1945 2694
rect 2001 2692 2025 2694
rect 2081 2692 2105 2694
rect 2161 2692 2185 2694
rect 2241 2692 2247 2694
rect 1939 2683 2247 2692
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2240 2446 2268 2586
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 2332 2310 2360 2790
rect 2424 2650 2452 3062
rect 2516 3058 2544 3334
rect 2599 3292 2907 3301
rect 2599 3290 2605 3292
rect 2661 3290 2685 3292
rect 2741 3290 2765 3292
rect 2821 3290 2845 3292
rect 2901 3290 2907 3292
rect 2661 3238 2663 3290
rect 2843 3238 2845 3290
rect 2599 3236 2605 3238
rect 2661 3236 2685 3238
rect 2741 3236 2765 3238
rect 2821 3236 2845 3238
rect 2901 3236 2907 3238
rect 2599 3227 2907 3236
rect 2976 3126 3004 3334
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2608 2582 2636 2858
rect 3068 2650 3096 3334
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2412 2508 2464 2514
rect 2464 2468 2544 2496
rect 2412 2450 2464 2456
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 1872 1970 1900 2246
rect 1860 1964 1912 1970
rect 1860 1906 1912 1912
rect 2516 1306 2544 2468
rect 2872 2440 2924 2446
rect 2924 2388 3004 2394
rect 2872 2382 3004 2388
rect 2884 2366 3004 2382
rect 2599 2204 2907 2213
rect 2599 2202 2605 2204
rect 2661 2202 2685 2204
rect 2741 2202 2765 2204
rect 2821 2202 2845 2204
rect 2901 2202 2907 2204
rect 2661 2150 2663 2202
rect 2843 2150 2845 2202
rect 2599 2148 2605 2150
rect 2661 2148 2685 2150
rect 2741 2148 2765 2150
rect 2821 2148 2845 2150
rect 2901 2148 2907 2150
rect 2599 2139 2907 2148
rect 2976 2038 3004 2366
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 2516 1278 2636 1306
rect 2608 800 2636 1278
rect 3252 800 3280 3470
rect 3344 2650 3372 3878
rect 3436 3194 3464 3998
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3528 2938 3556 3538
rect 3620 3398 3648 4014
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3436 2910 3556 2938
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 2446 3464 2910
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3528 2446 3556 2790
rect 3620 2446 3648 3130
rect 3712 2446 3740 4966
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 3618 3832 4422
rect 4172 4162 4200 4762
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4264 4282 4292 4626
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4172 4134 4292 4162
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3804 3590 3924 3618
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3804 1170 3832 3470
rect 3896 3466 3924 3590
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3896 3126 3924 3402
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3988 2854 4016 3674
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3126 4108 3538
rect 4160 3460 4212 3466
rect 4264 3448 4292 4134
rect 4356 4078 4384 4558
rect 4448 4282 4476 5188
rect 4620 5170 4672 5176
rect 4632 4826 4660 5170
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4816 4758 4844 5238
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4908 4554 4936 5358
rect 5092 5234 5120 5510
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4577 4380 4885 4389
rect 4577 4378 4583 4380
rect 4639 4378 4663 4380
rect 4719 4378 4743 4380
rect 4799 4378 4823 4380
rect 4879 4378 4885 4380
rect 4639 4326 4641 4378
rect 4821 4326 4823 4378
rect 4577 4324 4583 4326
rect 4639 4324 4663 4326
rect 4719 4324 4743 4326
rect 4799 4324 4823 4326
rect 4879 4324 4885 4326
rect 4577 4315 4885 4324
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4212 3420 4292 3448
rect 4448 3482 4476 4082
rect 5000 3602 5028 5102
rect 5092 4554 5120 5170
rect 5184 4690 5212 5850
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5368 5001 5396 5646
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5460 5098 5488 5578
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5354 4720 5410 4729
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 5184 4214 5212 4626
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4448 3466 4568 3482
rect 4448 3460 4580 3466
rect 4448 3454 4528 3460
rect 4160 3402 4212 3408
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4172 2922 4200 3402
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 3058 4384 3334
rect 4448 3194 4476 3454
rect 4528 3402 4580 3408
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4577 3292 4885 3301
rect 4577 3290 4583 3292
rect 4639 3290 4663 3292
rect 4719 3290 4743 3292
rect 4799 3290 4823 3292
rect 4879 3290 4885 3292
rect 4639 3238 4641 3290
rect 4821 3238 4823 3290
rect 4577 3236 4583 3238
rect 4639 3236 4663 3238
rect 4719 3236 4743 3238
rect 4799 3236 4823 3238
rect 4879 3236 4885 3238
rect 4577 3227 4885 3236
rect 5092 3194 5120 3334
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5184 3126 5212 4014
rect 5276 3738 5304 4694
rect 5354 4655 5410 4664
rect 5368 4146 5396 4655
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5552 4026 5580 5578
rect 5644 5370 5672 6190
rect 5736 5914 5764 6258
rect 6012 6100 6040 6598
rect 6288 6458 6316 7754
rect 6555 7644 6863 7653
rect 6555 7642 6561 7644
rect 6617 7642 6641 7644
rect 6697 7642 6721 7644
rect 6777 7642 6801 7644
rect 6857 7642 6863 7644
rect 6617 7590 6619 7642
rect 6799 7590 6801 7642
rect 6555 7588 6561 7590
rect 6617 7588 6641 7590
rect 6697 7588 6721 7590
rect 6777 7588 6801 7590
rect 6857 7588 6863 7590
rect 6555 7579 6863 7588
rect 6932 7528 6960 7890
rect 7024 7886 7052 8871
rect 7392 7954 7420 9318
rect 7576 9178 7604 9522
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8498 7604 9114
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7668 8634 7696 8910
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7760 8498 7788 9522
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7873 9276 8181 9285
rect 7873 9274 7879 9276
rect 7935 9274 7959 9276
rect 8015 9274 8039 9276
rect 8095 9274 8119 9276
rect 8175 9274 8181 9276
rect 7935 9222 7937 9274
rect 8117 9222 8119 9274
rect 7873 9220 7879 9222
rect 7935 9220 7959 9222
rect 8015 9220 8039 9222
rect 8095 9220 8119 9222
rect 8175 9220 8181 9222
rect 7873 9211 8181 9220
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7484 7954 7512 8230
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 6656 7500 6960 7528
rect 6656 7410 6684 7500
rect 6734 7440 6790 7449
rect 6644 7404 6696 7410
rect 7024 7410 7052 7686
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 6734 7375 6736 7384
rect 6644 7346 6696 7352
rect 6788 7375 6790 7384
rect 6920 7404 6972 7410
rect 6736 7346 6788 7352
rect 6920 7346 6972 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6932 6934 6960 7346
rect 7116 7002 7144 7346
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 5828 6072 6040 6100
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5828 5846 5856 6072
rect 5895 6012 6203 6021
rect 5895 6010 5901 6012
rect 5957 6010 5981 6012
rect 6037 6010 6061 6012
rect 6117 6010 6141 6012
rect 6197 6010 6203 6012
rect 5957 5958 5959 6010
rect 6139 5958 6141 6010
rect 5895 5956 5901 5958
rect 5957 5956 5981 5958
rect 6037 5956 6061 5958
rect 6117 5956 6141 5958
rect 6197 5956 6203 5958
rect 5895 5947 6203 5956
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5722 5264 5778 5273
rect 5632 5229 5684 5235
rect 5722 5199 5724 5208
rect 5632 5171 5684 5177
rect 5776 5199 5778 5208
rect 5644 4282 5672 5171
rect 5724 5170 5776 5176
rect 5828 4690 5856 5782
rect 5920 5642 5948 5850
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6012 5302 6040 5510
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5296 6052 5302
rect 6104 5273 6132 5306
rect 6000 5238 6052 5244
rect 6090 5264 6146 5273
rect 6196 5234 6224 5510
rect 6090 5199 6146 5208
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 5895 4924 6203 4933
rect 5895 4922 5901 4924
rect 5957 4922 5981 4924
rect 6037 4922 6061 4924
rect 6117 4922 6141 4924
rect 6197 4922 6203 4924
rect 5957 4870 5959 4922
rect 6139 4870 6141 4922
rect 5895 4868 5901 4870
rect 5957 4868 5981 4870
rect 6037 4868 6061 4870
rect 6117 4868 6141 4870
rect 6197 4868 6203 4870
rect 5895 4859 6203 4868
rect 6182 4720 6238 4729
rect 5816 4684 5868 4690
rect 6288 4690 6316 6190
rect 6380 6186 6408 6734
rect 6472 6304 6500 6870
rect 7208 6798 7236 7482
rect 7300 7002 7328 7686
rect 7484 7274 7512 7890
rect 7668 7750 7696 8230
rect 7760 8090 7788 8434
rect 8036 8430 8064 8978
rect 8208 8900 8260 8906
rect 8128 8860 8208 8888
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8128 8294 8156 8860
rect 8208 8842 8260 8848
rect 8312 8566 8340 9318
rect 8404 8974 8432 9386
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8300 8424 8352 8430
rect 8220 8372 8300 8378
rect 8220 8366 8352 8372
rect 8220 8350 8340 8366
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7873 8188 8181 8197
rect 7873 8186 7879 8188
rect 7935 8186 7959 8188
rect 8015 8186 8039 8188
rect 8095 8186 8119 8188
rect 8175 8186 8181 8188
rect 7935 8134 7937 8186
rect 8117 8134 8119 8186
rect 7873 8132 7879 8134
rect 7935 8132 7959 8134
rect 8015 8132 8039 8134
rect 8095 8132 8119 8134
rect 8175 8132 8181 8134
rect 7873 8123 8181 8132
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7760 7546 7788 7890
rect 8220 7886 8248 8350
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7852 7478 7880 7822
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7564 7336 7616 7342
rect 7562 7304 7564 7313
rect 7616 7304 7618 7313
rect 7472 7268 7524 7274
rect 7562 7239 7618 7248
rect 7472 7210 7524 7216
rect 7873 7100 8181 7109
rect 7873 7098 7879 7100
rect 7935 7098 7959 7100
rect 8015 7098 8039 7100
rect 8095 7098 8119 7100
rect 8175 7098 8181 7100
rect 7935 7046 7937 7098
rect 8117 7046 8119 7098
rect 7873 7044 7879 7046
rect 7935 7044 7959 7046
rect 8015 7044 8039 7046
rect 8095 7044 8119 7046
rect 8175 7044 8181 7046
rect 7873 7035 8181 7044
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6555 6556 6863 6565
rect 6555 6554 6561 6556
rect 6617 6554 6641 6556
rect 6697 6554 6721 6556
rect 6777 6554 6801 6556
rect 6857 6554 6863 6556
rect 6617 6502 6619 6554
rect 6799 6502 6801 6554
rect 6555 6500 6561 6502
rect 6617 6500 6641 6502
rect 6697 6500 6721 6502
rect 6777 6500 6801 6502
rect 6857 6500 6863 6502
rect 6555 6491 6863 6500
rect 6644 6452 6696 6458
rect 6696 6412 6868 6440
rect 6644 6394 6696 6400
rect 6552 6316 6604 6322
rect 6472 6276 6552 6304
rect 6552 6258 6604 6264
rect 6840 6202 6868 6412
rect 6932 6322 6960 6598
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6368 6180 6420 6186
rect 6840 6174 6960 6202
rect 6368 6122 6420 6128
rect 6368 5704 6420 5710
rect 6552 5704 6604 5710
rect 6368 5646 6420 5652
rect 6550 5672 6552 5681
rect 6604 5672 6606 5681
rect 6380 5234 6408 5646
rect 6932 5642 6960 6174
rect 7024 6118 7052 6598
rect 7116 6390 7144 6666
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7392 5914 7420 6734
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7484 5778 7512 6734
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 6550 5607 6606 5616
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6555 5468 6863 5477
rect 6555 5466 6561 5468
rect 6617 5466 6641 5468
rect 6697 5466 6721 5468
rect 6777 5466 6801 5468
rect 6857 5466 6863 5468
rect 6617 5414 6619 5466
rect 6799 5414 6801 5466
rect 6555 5412 6561 5414
rect 6617 5412 6641 5414
rect 6697 5412 6721 5414
rect 6777 5412 6801 5414
rect 6857 5412 6863 5414
rect 6555 5403 6863 5412
rect 6932 5352 6960 5578
rect 6840 5324 6960 5352
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6182 4655 6238 4664
rect 6276 4684 6328 4690
rect 5816 4626 5868 4632
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5368 3998 5580 4026
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5368 3602 5396 3998
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 4448 2650 4476 2858
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5276 2582 5304 3538
rect 5460 2582 5488 3878
rect 5552 3482 5580 3878
rect 5644 3738 5672 4082
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5736 3534 5764 4422
rect 6196 4146 6224 4655
rect 6276 4626 6328 4632
rect 6380 4146 6408 5170
rect 6748 4826 6776 5170
rect 6840 5166 6868 5324
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6840 4468 6868 5102
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6472 4440 6868 4468
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 5724 3528 5776 3534
rect 5552 3454 5672 3482
rect 5724 3470 5776 3476
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3058 5580 3334
rect 5644 3058 5672 3454
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5552 2514 5580 2586
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4068 2304 4120 2310
rect 4172 2292 4200 2382
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 4120 2264 4200 2292
rect 4068 2246 4120 2252
rect 4448 1170 4476 2314
rect 4577 2204 4885 2213
rect 4577 2202 4583 2204
rect 4639 2202 4663 2204
rect 4719 2202 4743 2204
rect 4799 2202 4823 2204
rect 4879 2202 4885 2204
rect 4639 2150 4641 2202
rect 4821 2150 4823 2202
rect 4577 2148 4583 2150
rect 4639 2148 4663 2150
rect 4719 2148 4743 2150
rect 4799 2148 4823 2150
rect 4879 2148 4885 2150
rect 4577 2139 4885 2148
rect 3804 1142 3924 1170
rect 4448 1142 4568 1170
rect 3896 800 3924 1142
rect 4540 800 4568 1142
rect 5184 800 5212 2314
rect 5552 1970 5580 2450
rect 5736 2446 5764 2790
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5828 2310 5856 4082
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 5895 3836 6203 3845
rect 5895 3834 5901 3836
rect 5957 3834 5981 3836
rect 6037 3834 6061 3836
rect 6117 3834 6141 3836
rect 6197 3834 6203 3836
rect 5957 3782 5959 3834
rect 6139 3782 6141 3834
rect 5895 3780 5901 3782
rect 5957 3780 5981 3782
rect 6037 3780 6061 3782
rect 6117 3780 6141 3782
rect 6197 3780 6203 3782
rect 5895 3771 6203 3780
rect 5895 2748 6203 2757
rect 5895 2746 5901 2748
rect 5957 2746 5981 2748
rect 6037 2746 6061 2748
rect 6117 2746 6141 2748
rect 6197 2746 6203 2748
rect 5957 2694 5959 2746
rect 6139 2694 6141 2746
rect 5895 2692 5901 2694
rect 5957 2692 5981 2694
rect 6037 2692 6061 2694
rect 6117 2692 6141 2694
rect 6197 2692 6203 2694
rect 5895 2683 6203 2692
rect 6288 2650 6316 4014
rect 6380 4010 6408 4082
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 2650 6408 3402
rect 6472 3176 6500 4440
rect 6555 4380 6863 4389
rect 6555 4378 6561 4380
rect 6617 4378 6641 4380
rect 6697 4378 6721 4380
rect 6777 4378 6801 4380
rect 6857 4378 6863 4380
rect 6617 4326 6619 4378
rect 6799 4326 6801 4378
rect 6555 4324 6561 4326
rect 6617 4324 6641 4326
rect 6697 4324 6721 4326
rect 6777 4324 6801 4326
rect 6857 4324 6863 4326
rect 6555 4315 6863 4324
rect 6932 4078 6960 5034
rect 7116 4282 7144 5646
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 4690 7236 5510
rect 7392 5098 7420 5646
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7010 4176 7066 4185
rect 7010 4111 7066 4120
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6932 3754 6960 4014
rect 6840 3726 6960 3754
rect 6840 3398 6868 3726
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6555 3292 6863 3301
rect 6555 3290 6561 3292
rect 6617 3290 6641 3292
rect 6697 3290 6721 3292
rect 6777 3290 6801 3292
rect 6857 3290 6863 3292
rect 6617 3238 6619 3290
rect 6799 3238 6801 3290
rect 6555 3236 6561 3238
rect 6617 3236 6641 3238
rect 6697 3236 6721 3238
rect 6777 3236 6801 3238
rect 6857 3236 6863 3238
rect 6555 3227 6863 3236
rect 6644 3188 6696 3194
rect 6472 3148 6592 3176
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6288 2310 6316 2586
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6000 2032 6052 2038
rect 5998 2000 6000 2009
rect 6052 2000 6054 2009
rect 5540 1964 5592 1970
rect 5998 1935 6054 1944
rect 5540 1906 5592 1912
rect 6472 800 6500 2790
rect 6564 2446 6592 3148
rect 6644 3130 6696 3136
rect 6656 3058 6684 3130
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6840 2378 6868 2926
rect 6932 2446 6960 3606
rect 7024 3534 7052 4111
rect 7116 4078 7144 4218
rect 7208 4214 7236 4626
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7300 4146 7328 5034
rect 7392 4146 7420 5034
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7300 3670 7328 4082
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7208 3074 7236 3470
rect 7484 3194 7512 5578
rect 7576 4282 7604 6666
rect 8128 6458 8156 6734
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7668 4690 7696 6054
rect 7760 5778 7788 6054
rect 7873 6012 8181 6021
rect 7873 6010 7879 6012
rect 7935 6010 7959 6012
rect 8015 6010 8039 6012
rect 8095 6010 8119 6012
rect 8175 6010 8181 6012
rect 7935 5958 7937 6010
rect 8117 5958 8119 6010
rect 7873 5956 7879 5958
rect 7935 5956 7959 5958
rect 8015 5956 8039 5958
rect 8095 5956 8119 5958
rect 8175 5956 8181 5958
rect 7873 5947 8181 5956
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7944 5710 7972 5782
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8024 5704 8076 5710
rect 8220 5692 8248 7686
rect 8312 7410 8340 7822
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8404 7290 8432 8774
rect 8533 8732 8841 8741
rect 8533 8730 8539 8732
rect 8595 8730 8619 8732
rect 8675 8730 8699 8732
rect 8755 8730 8779 8732
rect 8835 8730 8841 8732
rect 8595 8678 8597 8730
rect 8777 8678 8779 8730
rect 8533 8676 8539 8678
rect 8595 8676 8619 8678
rect 8675 8676 8699 8678
rect 8755 8676 8779 8678
rect 8835 8676 8841 8678
rect 8533 8667 8841 8676
rect 8956 8265 8984 9522
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 8430 9076 8842
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8942 8256 8998 8265
rect 8942 8191 8998 8200
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8533 7644 8841 7653
rect 8533 7642 8539 7644
rect 8595 7642 8619 7644
rect 8675 7642 8699 7644
rect 8755 7642 8779 7644
rect 8835 7642 8841 7644
rect 8595 7590 8597 7642
rect 8777 7590 8779 7642
rect 8533 7588 8539 7590
rect 8595 7588 8619 7590
rect 8675 7588 8699 7590
rect 8755 7588 8779 7590
rect 8835 7588 8841 7590
rect 8533 7579 8841 7588
rect 8956 7585 8984 7686
rect 8942 7576 8998 7585
rect 8942 7511 8998 7520
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8076 5664 8248 5692
rect 8312 7262 8432 7290
rect 8024 5646 8076 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7873 4924 8181 4933
rect 7873 4922 7879 4924
rect 7935 4922 7959 4924
rect 8015 4922 8039 4924
rect 8095 4922 8119 4924
rect 8175 4922 8181 4924
rect 7935 4870 7937 4922
rect 8117 4870 8119 4922
rect 7873 4868 7879 4870
rect 7935 4868 7959 4870
rect 8015 4868 8039 4870
rect 8095 4868 8119 4870
rect 8175 4868 8181 4870
rect 7873 4859 8181 4868
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7668 4078 7696 4626
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7760 3602 7788 4558
rect 8220 4146 8248 5510
rect 8312 4826 8340 7262
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 5642 8432 7142
rect 8496 6662 8524 7346
rect 8588 6905 8616 7346
rect 8574 6896 8630 6905
rect 8574 6831 8630 6840
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8533 6556 8841 6565
rect 8533 6554 8539 6556
rect 8595 6554 8619 6556
rect 8675 6554 8699 6556
rect 8755 6554 8779 6556
rect 8835 6554 8841 6556
rect 8595 6502 8597 6554
rect 8777 6502 8779 6554
rect 8533 6500 8539 6502
rect 8595 6500 8619 6502
rect 8675 6500 8699 6502
rect 8755 6500 8779 6502
rect 8835 6500 8841 6502
rect 8533 6491 8841 6500
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8496 5574 8524 6394
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8588 6225 8616 6258
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8956 5846 8984 6666
rect 9048 6458 9076 8366
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9140 7449 9168 8298
rect 9126 7440 9182 7449
rect 9126 7375 9182 7384
rect 9140 6730 9168 7375
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8942 5536 8998 5545
rect 8533 5468 8841 5477
rect 8942 5471 8998 5480
rect 8533 5466 8539 5468
rect 8595 5466 8619 5468
rect 8675 5466 8699 5468
rect 8755 5466 8779 5468
rect 8835 5466 8841 5468
rect 8595 5414 8597 5466
rect 8777 5414 8779 5466
rect 8533 5412 8539 5414
rect 8595 5412 8619 5414
rect 8675 5412 8699 5414
rect 8755 5412 8779 5414
rect 8835 5412 8841 5414
rect 8533 5403 8841 5412
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8404 4146 8432 4966
rect 8533 4380 8841 4389
rect 8533 4378 8539 4380
rect 8595 4378 8619 4380
rect 8675 4378 8699 4380
rect 8755 4378 8779 4380
rect 8835 4378 8841 4380
rect 8595 4326 8597 4378
rect 8777 4326 8779 4378
rect 8533 4324 8539 4326
rect 8595 4324 8619 4326
rect 8675 4324 8699 4326
rect 8755 4324 8779 4326
rect 8835 4324 8841 4326
rect 8533 4315 8841 4324
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 7873 3836 8181 3845
rect 7873 3834 7879 3836
rect 7935 3834 7959 3836
rect 8015 3834 8039 3836
rect 8095 3834 8119 3836
rect 8175 3834 8181 3836
rect 7935 3782 7937 3834
rect 8117 3782 8119 3834
rect 7873 3780 7879 3782
rect 7935 3780 7959 3782
rect 8015 3780 8039 3782
rect 8095 3780 8119 3782
rect 8175 3780 8181 3782
rect 7873 3771 8181 3780
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7208 3046 7328 3074
rect 7392 3058 7420 3130
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7024 2650 7052 2926
rect 7300 2854 7328 3046
rect 7380 3052 7432 3058
rect 7432 3012 7512 3040
rect 7380 2994 7432 3000
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7378 2816 7434 2825
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7208 2446 7236 2790
rect 7300 2446 7328 2790
rect 7378 2751 7434 2760
rect 7392 2650 7420 2751
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2514 7512 3012
rect 7576 2650 7604 3470
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7760 3058 7788 3402
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7852 2990 7880 3130
rect 8128 3058 8156 3334
rect 8220 3058 8248 3606
rect 8312 3194 8340 4082
rect 8956 4010 8984 5471
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8496 3505 8524 3674
rect 8482 3496 8538 3505
rect 8392 3460 8444 3466
rect 8482 3431 8538 3440
rect 8392 3402 8444 3408
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7760 2825 7788 2858
rect 8300 2848 8352 2854
rect 7746 2816 7802 2825
rect 8300 2790 8352 2796
rect 7746 2751 7802 2760
rect 7873 2748 8181 2757
rect 7873 2746 7879 2748
rect 7935 2746 7959 2748
rect 8015 2746 8039 2748
rect 8095 2746 8119 2748
rect 8175 2746 8181 2748
rect 7935 2694 7937 2746
rect 8117 2694 8119 2746
rect 7873 2692 7879 2694
rect 7935 2692 7959 2694
rect 8015 2692 8039 2694
rect 8095 2692 8119 2694
rect 8175 2692 8181 2694
rect 7873 2683 8181 2692
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 8312 2446 8340 2790
rect 8404 2650 8432 3402
rect 8533 3292 8841 3301
rect 8533 3290 8539 3292
rect 8595 3290 8619 3292
rect 8675 3290 8699 3292
rect 8755 3290 8779 3292
rect 8835 3290 8841 3292
rect 8595 3238 8597 3290
rect 8777 3238 8779 3290
rect 8533 3236 8539 3238
rect 8595 3236 8619 3238
rect 8675 3236 8699 3238
rect 8755 3236 8779 3238
rect 8835 3236 8841 3238
rect 8533 3227 8841 3236
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6555 2204 6863 2213
rect 6555 2202 6561 2204
rect 6617 2202 6641 2204
rect 6697 2202 6721 2204
rect 6777 2202 6801 2204
rect 6857 2202 6863 2204
rect 6617 2150 6619 2202
rect 6799 2150 6801 2202
rect 6555 2148 6561 2150
rect 6617 2148 6641 2150
rect 6697 2148 6721 2150
rect 6777 2148 6801 2150
rect 6857 2148 6863 2150
rect 6555 2139 6863 2148
rect 8533 2204 8841 2213
rect 8533 2202 8539 2204
rect 8595 2202 8619 2204
rect 8675 2202 8699 2204
rect 8755 2202 8779 2204
rect 8835 2202 8841 2204
rect 8595 2150 8597 2202
rect 8777 2150 8779 2202
rect 8533 2148 8539 2150
rect 8595 2148 8619 2150
rect 8675 2148 8699 2150
rect 8755 2148 8779 2150
rect 8835 2148 8841 2150
rect 8533 2139 8841 2148
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
<< via2 >>
rect 2605 9818 2661 9820
rect 2685 9818 2741 9820
rect 2765 9818 2821 9820
rect 2845 9818 2901 9820
rect 2605 9766 2651 9818
rect 2651 9766 2661 9818
rect 2685 9766 2715 9818
rect 2715 9766 2727 9818
rect 2727 9766 2741 9818
rect 2765 9766 2779 9818
rect 2779 9766 2791 9818
rect 2791 9766 2821 9818
rect 2845 9766 2855 9818
rect 2855 9766 2901 9818
rect 2605 9764 2661 9766
rect 2685 9764 2741 9766
rect 2765 9764 2821 9766
rect 2845 9764 2901 9766
rect 4583 9818 4639 9820
rect 4663 9818 4719 9820
rect 4743 9818 4799 9820
rect 4823 9818 4879 9820
rect 4583 9766 4629 9818
rect 4629 9766 4639 9818
rect 4663 9766 4693 9818
rect 4693 9766 4705 9818
rect 4705 9766 4719 9818
rect 4743 9766 4757 9818
rect 4757 9766 4769 9818
rect 4769 9766 4799 9818
rect 4823 9766 4833 9818
rect 4833 9766 4879 9818
rect 4583 9764 4639 9766
rect 4663 9764 4719 9766
rect 4743 9764 4799 9766
rect 4823 9764 4879 9766
rect 6561 9818 6617 9820
rect 6641 9818 6697 9820
rect 6721 9818 6777 9820
rect 6801 9818 6857 9820
rect 6561 9766 6607 9818
rect 6607 9766 6617 9818
rect 6641 9766 6671 9818
rect 6671 9766 6683 9818
rect 6683 9766 6697 9818
rect 6721 9766 6735 9818
rect 6735 9766 6747 9818
rect 6747 9766 6777 9818
rect 6801 9766 6811 9818
rect 6811 9766 6857 9818
rect 6561 9764 6617 9766
rect 6641 9764 6697 9766
rect 6721 9764 6777 9766
rect 6801 9764 6857 9766
rect 8539 9818 8595 9820
rect 8619 9818 8675 9820
rect 8699 9818 8755 9820
rect 8779 9818 8835 9820
rect 8539 9766 8585 9818
rect 8585 9766 8595 9818
rect 8619 9766 8649 9818
rect 8649 9766 8661 9818
rect 8661 9766 8675 9818
rect 8699 9766 8713 9818
rect 8713 9766 8725 9818
rect 8725 9766 8755 9818
rect 8779 9766 8789 9818
rect 8789 9766 8835 9818
rect 8539 9764 8595 9766
rect 8619 9764 8675 9766
rect 8699 9764 8755 9766
rect 8779 9764 8835 9766
rect 1030 9596 1032 9616
rect 1032 9596 1084 9616
rect 1084 9596 1086 9616
rect 1030 9560 1086 9596
rect 1398 8880 1454 8936
rect 1945 9274 2001 9276
rect 2025 9274 2081 9276
rect 2105 9274 2161 9276
rect 2185 9274 2241 9276
rect 1945 9222 1991 9274
rect 1991 9222 2001 9274
rect 2025 9222 2055 9274
rect 2055 9222 2067 9274
rect 2067 9222 2081 9274
rect 2105 9222 2119 9274
rect 2119 9222 2131 9274
rect 2131 9222 2161 9274
rect 2185 9222 2195 9274
rect 2195 9222 2241 9274
rect 1945 9220 2001 9222
rect 2025 9220 2081 9222
rect 2105 9220 2161 9222
rect 2185 9220 2241 9222
rect 1490 8200 1546 8256
rect 1306 7520 1362 7576
rect 846 6604 848 6624
rect 848 6604 900 6624
rect 900 6604 902 6624
rect 846 6568 902 6604
rect 1945 8186 2001 8188
rect 2025 8186 2081 8188
rect 2105 8186 2161 8188
rect 2185 8186 2241 8188
rect 1945 8134 1991 8186
rect 1991 8134 2001 8186
rect 2025 8134 2055 8186
rect 2055 8134 2067 8186
rect 2067 8134 2081 8186
rect 2105 8134 2119 8186
rect 2119 8134 2131 8186
rect 2131 8134 2161 8186
rect 2185 8134 2195 8186
rect 2195 8134 2241 8186
rect 1945 8132 2001 8134
rect 2025 8132 2081 8134
rect 2105 8132 2161 8134
rect 2185 8132 2241 8134
rect 846 5888 902 5944
rect 1398 5752 1454 5808
rect 938 5480 994 5536
rect 2605 8730 2661 8732
rect 2685 8730 2741 8732
rect 2765 8730 2821 8732
rect 2845 8730 2901 8732
rect 2605 8678 2651 8730
rect 2651 8678 2661 8730
rect 2685 8678 2715 8730
rect 2715 8678 2727 8730
rect 2727 8678 2741 8730
rect 2765 8678 2779 8730
rect 2779 8678 2791 8730
rect 2791 8678 2821 8730
rect 2845 8678 2855 8730
rect 2855 8678 2901 8730
rect 2605 8676 2661 8678
rect 2685 8676 2741 8678
rect 2765 8676 2821 8678
rect 2845 8676 2901 8678
rect 3923 9274 3979 9276
rect 4003 9274 4059 9276
rect 4083 9274 4139 9276
rect 4163 9274 4219 9276
rect 3923 9222 3969 9274
rect 3969 9222 3979 9274
rect 4003 9222 4033 9274
rect 4033 9222 4045 9274
rect 4045 9222 4059 9274
rect 4083 9222 4097 9274
rect 4097 9222 4109 9274
rect 4109 9222 4139 9274
rect 4163 9222 4173 9274
rect 4173 9222 4219 9274
rect 3923 9220 3979 9222
rect 4003 9220 4059 9222
rect 4083 9220 4139 9222
rect 4163 9220 4219 9222
rect 1945 7098 2001 7100
rect 2025 7098 2081 7100
rect 2105 7098 2161 7100
rect 2185 7098 2241 7100
rect 1945 7046 1991 7098
rect 1991 7046 2001 7098
rect 2025 7046 2055 7098
rect 2055 7046 2067 7098
rect 2067 7046 2081 7098
rect 2105 7046 2119 7098
rect 2119 7046 2131 7098
rect 2131 7046 2161 7098
rect 2185 7046 2195 7098
rect 2195 7046 2241 7098
rect 1945 7044 2001 7046
rect 2025 7044 2081 7046
rect 2105 7044 2161 7046
rect 2185 7044 2241 7046
rect 1945 6010 2001 6012
rect 2025 6010 2081 6012
rect 2105 6010 2161 6012
rect 2185 6010 2241 6012
rect 1945 5958 1991 6010
rect 1991 5958 2001 6010
rect 2025 5958 2055 6010
rect 2055 5958 2067 6010
rect 2067 5958 2081 6010
rect 2105 5958 2119 6010
rect 2119 5958 2131 6010
rect 2131 5958 2161 6010
rect 2185 5958 2195 6010
rect 2195 5958 2241 6010
rect 1945 5956 2001 5958
rect 2025 5956 2081 5958
rect 2105 5956 2161 5958
rect 2185 5956 2241 5958
rect 2605 7642 2661 7644
rect 2685 7642 2741 7644
rect 2765 7642 2821 7644
rect 2845 7642 2901 7644
rect 2605 7590 2651 7642
rect 2651 7590 2661 7642
rect 2685 7590 2715 7642
rect 2715 7590 2727 7642
rect 2727 7590 2741 7642
rect 2765 7590 2779 7642
rect 2779 7590 2791 7642
rect 2791 7590 2821 7642
rect 2845 7590 2855 7642
rect 2855 7590 2901 7642
rect 2605 7588 2661 7590
rect 2685 7588 2741 7590
rect 2765 7588 2821 7590
rect 2845 7588 2901 7590
rect 2605 6554 2661 6556
rect 2685 6554 2741 6556
rect 2765 6554 2821 6556
rect 2845 6554 2901 6556
rect 2605 6502 2651 6554
rect 2651 6502 2661 6554
rect 2685 6502 2715 6554
rect 2715 6502 2727 6554
rect 2727 6502 2741 6554
rect 2765 6502 2779 6554
rect 2779 6502 2791 6554
rect 2791 6502 2821 6554
rect 2845 6502 2855 6554
rect 2855 6502 2901 6554
rect 2605 6500 2661 6502
rect 2685 6500 2741 6502
rect 2765 6500 2821 6502
rect 2845 6500 2901 6502
rect 1490 4800 1546 4856
rect 1945 4922 2001 4924
rect 2025 4922 2081 4924
rect 2105 4922 2161 4924
rect 2185 4922 2241 4924
rect 1945 4870 1991 4922
rect 1991 4870 2001 4922
rect 2025 4870 2055 4922
rect 2055 4870 2067 4922
rect 2067 4870 2081 4922
rect 2105 4870 2119 4922
rect 2119 4870 2131 4922
rect 2131 4870 2161 4922
rect 2185 4870 2195 4922
rect 2195 4870 2241 4922
rect 1945 4868 2001 4870
rect 2025 4868 2081 4870
rect 2105 4868 2161 4870
rect 2185 4868 2241 4870
rect 2605 5466 2661 5468
rect 2685 5466 2741 5468
rect 2765 5466 2821 5468
rect 2845 5466 2901 5468
rect 2605 5414 2651 5466
rect 2651 5414 2661 5466
rect 2685 5414 2715 5466
rect 2715 5414 2727 5466
rect 2727 5414 2741 5466
rect 2765 5414 2779 5466
rect 2779 5414 2791 5466
rect 2791 5414 2821 5466
rect 2845 5414 2855 5466
rect 2855 5414 2901 5466
rect 2605 5412 2661 5414
rect 2685 5412 2741 5414
rect 2765 5412 2821 5414
rect 2845 5412 2901 5414
rect 2605 4378 2661 4380
rect 2685 4378 2741 4380
rect 2765 4378 2821 4380
rect 2845 4378 2901 4380
rect 2605 4326 2651 4378
rect 2651 4326 2661 4378
rect 2685 4326 2715 4378
rect 2715 4326 2727 4378
rect 2727 4326 2741 4378
rect 2765 4326 2779 4378
rect 2779 4326 2791 4378
rect 2791 4326 2821 4378
rect 2845 4326 2855 4378
rect 2855 4326 2901 4378
rect 2605 4324 2661 4326
rect 2685 4324 2741 4326
rect 2765 4324 2821 4326
rect 2845 4324 2901 4326
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 1945 3834 2001 3836
rect 2025 3834 2081 3836
rect 2105 3834 2161 3836
rect 2185 3834 2241 3836
rect 1945 3782 1991 3834
rect 1991 3782 2001 3834
rect 2025 3782 2055 3834
rect 2055 3782 2067 3834
rect 2067 3782 2081 3834
rect 2105 3782 2119 3834
rect 2119 3782 2131 3834
rect 2131 3782 2161 3834
rect 2185 3782 2195 3834
rect 2195 3782 2241 3834
rect 1945 3780 2001 3782
rect 2025 3780 2081 3782
rect 2105 3780 2161 3782
rect 2185 3780 2241 3782
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 4583 8730 4639 8732
rect 4663 8730 4719 8732
rect 4743 8730 4799 8732
rect 4823 8730 4879 8732
rect 4583 8678 4629 8730
rect 4629 8678 4639 8730
rect 4663 8678 4693 8730
rect 4693 8678 4705 8730
rect 4705 8678 4719 8730
rect 4743 8678 4757 8730
rect 4757 8678 4769 8730
rect 4769 8678 4799 8730
rect 4823 8678 4833 8730
rect 4833 8678 4879 8730
rect 4583 8676 4639 8678
rect 4663 8676 4719 8678
rect 4743 8676 4799 8678
rect 4823 8676 4879 8678
rect 4583 7642 4639 7644
rect 4663 7642 4719 7644
rect 4743 7642 4799 7644
rect 4823 7642 4879 7644
rect 4583 7590 4629 7642
rect 4629 7590 4639 7642
rect 4663 7590 4693 7642
rect 4693 7590 4705 7642
rect 4705 7590 4719 7642
rect 4743 7590 4757 7642
rect 4757 7590 4769 7642
rect 4769 7590 4799 7642
rect 4823 7590 4833 7642
rect 4833 7590 4879 7642
rect 4583 7588 4639 7590
rect 4663 7588 4719 7590
rect 4743 7588 4799 7590
rect 4823 7588 4879 7590
rect 5901 9274 5957 9276
rect 5981 9274 6037 9276
rect 6061 9274 6117 9276
rect 6141 9274 6197 9276
rect 5901 9222 5947 9274
rect 5947 9222 5957 9274
rect 5981 9222 6011 9274
rect 6011 9222 6023 9274
rect 6023 9222 6037 9274
rect 6061 9222 6075 9274
rect 6075 9222 6087 9274
rect 6087 9222 6117 9274
rect 6141 9222 6151 9274
rect 6151 9222 6197 9274
rect 5901 9220 5957 9222
rect 5981 9220 6037 9222
rect 6061 9220 6117 9222
rect 6141 9220 6197 9222
rect 7010 8880 7066 8936
rect 6561 8730 6617 8732
rect 6641 8730 6697 8732
rect 6721 8730 6777 8732
rect 6801 8730 6857 8732
rect 6561 8678 6607 8730
rect 6607 8678 6617 8730
rect 6641 8678 6671 8730
rect 6671 8678 6683 8730
rect 6683 8678 6697 8730
rect 6721 8678 6735 8730
rect 6735 8678 6747 8730
rect 6747 8678 6777 8730
rect 6801 8678 6811 8730
rect 6811 8678 6857 8730
rect 6561 8676 6617 8678
rect 6641 8676 6697 8678
rect 6721 8676 6777 8678
rect 6801 8676 6857 8678
rect 5901 8186 5957 8188
rect 5981 8186 6037 8188
rect 6061 8186 6117 8188
rect 6141 8186 6197 8188
rect 5901 8134 5947 8186
rect 5947 8134 5957 8186
rect 5981 8134 6011 8186
rect 6011 8134 6023 8186
rect 6023 8134 6037 8186
rect 6061 8134 6075 8186
rect 6075 8134 6087 8186
rect 6087 8134 6117 8186
rect 6141 8134 6151 8186
rect 6151 8134 6197 8186
rect 5901 8132 5957 8134
rect 5981 8132 6037 8134
rect 6061 8132 6117 8134
rect 6141 8132 6197 8134
rect 4583 6554 4639 6556
rect 4663 6554 4719 6556
rect 4743 6554 4799 6556
rect 4823 6554 4879 6556
rect 4583 6502 4629 6554
rect 4629 6502 4639 6554
rect 4663 6502 4693 6554
rect 4693 6502 4705 6554
rect 4705 6502 4719 6554
rect 4743 6502 4757 6554
rect 4757 6502 4769 6554
rect 4769 6502 4799 6554
rect 4823 6502 4833 6554
rect 4833 6502 4879 6554
rect 4583 6500 4639 6502
rect 4663 6500 4719 6502
rect 4743 6500 4799 6502
rect 4823 6500 4879 6502
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 4342 5772 4398 5808
rect 5354 7248 5410 7304
rect 5901 7098 5957 7100
rect 5981 7098 6037 7100
rect 6061 7098 6117 7100
rect 6141 7098 6197 7100
rect 5901 7046 5947 7098
rect 5947 7046 5957 7098
rect 5981 7046 6011 7098
rect 6011 7046 6023 7098
rect 6023 7046 6037 7098
rect 6061 7046 6075 7098
rect 6075 7046 6087 7098
rect 6087 7046 6117 7098
rect 6141 7046 6151 7098
rect 6151 7046 6197 7098
rect 5901 7044 5957 7046
rect 5981 7044 6037 7046
rect 6061 7044 6117 7046
rect 6141 7044 6197 7046
rect 4342 5752 4344 5772
rect 4344 5752 4396 5772
rect 4396 5752 4398 5772
rect 4583 5466 4639 5468
rect 4663 5466 4719 5468
rect 4743 5466 4799 5468
rect 4823 5466 4879 5468
rect 4583 5414 4629 5466
rect 4629 5414 4639 5466
rect 4663 5414 4693 5466
rect 4693 5414 4705 5466
rect 4705 5414 4719 5466
rect 4743 5414 4757 5466
rect 4757 5414 4769 5466
rect 4769 5414 4799 5466
rect 4823 5414 4833 5466
rect 4833 5414 4879 5466
rect 4583 5412 4639 5414
rect 4663 5412 4719 5414
rect 4743 5412 4799 5414
rect 4823 5412 4879 5414
rect 5078 5616 5134 5672
rect 1945 2746 2001 2748
rect 2025 2746 2081 2748
rect 2105 2746 2161 2748
rect 2185 2746 2241 2748
rect 1674 2488 1730 2544
rect 1945 2694 1991 2746
rect 1991 2694 2001 2746
rect 2025 2694 2055 2746
rect 2055 2694 2067 2746
rect 2067 2694 2081 2746
rect 2105 2694 2119 2746
rect 2119 2694 2131 2746
rect 2131 2694 2161 2746
rect 2185 2694 2195 2746
rect 2195 2694 2241 2746
rect 1945 2692 2001 2694
rect 2025 2692 2081 2694
rect 2105 2692 2161 2694
rect 2185 2692 2241 2694
rect 2605 3290 2661 3292
rect 2685 3290 2741 3292
rect 2765 3290 2821 3292
rect 2845 3290 2901 3292
rect 2605 3238 2651 3290
rect 2651 3238 2661 3290
rect 2685 3238 2715 3290
rect 2715 3238 2727 3290
rect 2727 3238 2741 3290
rect 2765 3238 2779 3290
rect 2779 3238 2791 3290
rect 2791 3238 2821 3290
rect 2845 3238 2855 3290
rect 2855 3238 2901 3290
rect 2605 3236 2661 3238
rect 2685 3236 2741 3238
rect 2765 3236 2821 3238
rect 2845 3236 2901 3238
rect 2605 2202 2661 2204
rect 2685 2202 2741 2204
rect 2765 2202 2821 2204
rect 2845 2202 2901 2204
rect 2605 2150 2651 2202
rect 2651 2150 2661 2202
rect 2685 2150 2715 2202
rect 2715 2150 2727 2202
rect 2727 2150 2741 2202
rect 2765 2150 2779 2202
rect 2779 2150 2791 2202
rect 2791 2150 2821 2202
rect 2845 2150 2855 2202
rect 2855 2150 2901 2202
rect 2605 2148 2661 2150
rect 2685 2148 2741 2150
rect 2765 2148 2821 2150
rect 2845 2148 2901 2150
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 4583 4378 4639 4380
rect 4663 4378 4719 4380
rect 4743 4378 4799 4380
rect 4823 4378 4879 4380
rect 4583 4326 4629 4378
rect 4629 4326 4639 4378
rect 4663 4326 4693 4378
rect 4693 4326 4705 4378
rect 4705 4326 4719 4378
rect 4743 4326 4757 4378
rect 4757 4326 4769 4378
rect 4769 4326 4799 4378
rect 4823 4326 4833 4378
rect 4833 4326 4879 4378
rect 4583 4324 4639 4326
rect 4663 4324 4719 4326
rect 4743 4324 4799 4326
rect 4823 4324 4879 4326
rect 5354 4936 5410 4992
rect 4583 3290 4639 3292
rect 4663 3290 4719 3292
rect 4743 3290 4799 3292
rect 4823 3290 4879 3292
rect 4583 3238 4629 3290
rect 4629 3238 4639 3290
rect 4663 3238 4693 3290
rect 4693 3238 4705 3290
rect 4705 3238 4719 3290
rect 4743 3238 4757 3290
rect 4757 3238 4769 3290
rect 4769 3238 4799 3290
rect 4823 3238 4833 3290
rect 4833 3238 4879 3290
rect 4583 3236 4639 3238
rect 4663 3236 4719 3238
rect 4743 3236 4799 3238
rect 4823 3236 4879 3238
rect 5354 4664 5410 4720
rect 6561 7642 6617 7644
rect 6641 7642 6697 7644
rect 6721 7642 6777 7644
rect 6801 7642 6857 7644
rect 6561 7590 6607 7642
rect 6607 7590 6617 7642
rect 6641 7590 6671 7642
rect 6671 7590 6683 7642
rect 6683 7590 6697 7642
rect 6721 7590 6735 7642
rect 6735 7590 6747 7642
rect 6747 7590 6777 7642
rect 6801 7590 6811 7642
rect 6811 7590 6857 7642
rect 6561 7588 6617 7590
rect 6641 7588 6697 7590
rect 6721 7588 6777 7590
rect 6801 7588 6857 7590
rect 7879 9274 7935 9276
rect 7959 9274 8015 9276
rect 8039 9274 8095 9276
rect 8119 9274 8175 9276
rect 7879 9222 7925 9274
rect 7925 9222 7935 9274
rect 7959 9222 7989 9274
rect 7989 9222 8001 9274
rect 8001 9222 8015 9274
rect 8039 9222 8053 9274
rect 8053 9222 8065 9274
rect 8065 9222 8095 9274
rect 8119 9222 8129 9274
rect 8129 9222 8175 9274
rect 7879 9220 7935 9222
rect 7959 9220 8015 9222
rect 8039 9220 8095 9222
rect 8119 9220 8175 9222
rect 6734 7404 6790 7440
rect 6734 7384 6736 7404
rect 6736 7384 6788 7404
rect 6788 7384 6790 7404
rect 5901 6010 5957 6012
rect 5981 6010 6037 6012
rect 6061 6010 6117 6012
rect 6141 6010 6197 6012
rect 5901 5958 5947 6010
rect 5947 5958 5957 6010
rect 5981 5958 6011 6010
rect 6011 5958 6023 6010
rect 6023 5958 6037 6010
rect 6061 5958 6075 6010
rect 6075 5958 6087 6010
rect 6087 5958 6117 6010
rect 6141 5958 6151 6010
rect 6151 5958 6197 6010
rect 5901 5956 5957 5958
rect 5981 5956 6037 5958
rect 6061 5956 6117 5958
rect 6141 5956 6197 5958
rect 5722 5228 5778 5264
rect 5722 5208 5724 5228
rect 5724 5208 5776 5228
rect 5776 5208 5778 5228
rect 6090 5208 6146 5264
rect 5901 4922 5957 4924
rect 5981 4922 6037 4924
rect 6061 4922 6117 4924
rect 6141 4922 6197 4924
rect 5901 4870 5947 4922
rect 5947 4870 5957 4922
rect 5981 4870 6011 4922
rect 6011 4870 6023 4922
rect 6023 4870 6037 4922
rect 6061 4870 6075 4922
rect 6075 4870 6087 4922
rect 6087 4870 6117 4922
rect 6141 4870 6151 4922
rect 6151 4870 6197 4922
rect 5901 4868 5957 4870
rect 5981 4868 6037 4870
rect 6061 4868 6117 4870
rect 6141 4868 6197 4870
rect 6182 4664 6238 4720
rect 7879 8186 7935 8188
rect 7959 8186 8015 8188
rect 8039 8186 8095 8188
rect 8119 8186 8175 8188
rect 7879 8134 7925 8186
rect 7925 8134 7935 8186
rect 7959 8134 7989 8186
rect 7989 8134 8001 8186
rect 8001 8134 8015 8186
rect 8039 8134 8053 8186
rect 8053 8134 8065 8186
rect 8065 8134 8095 8186
rect 8119 8134 8129 8186
rect 8129 8134 8175 8186
rect 7879 8132 7935 8134
rect 7959 8132 8015 8134
rect 8039 8132 8095 8134
rect 8119 8132 8175 8134
rect 7562 7284 7564 7304
rect 7564 7284 7616 7304
rect 7616 7284 7618 7304
rect 7562 7248 7618 7284
rect 7879 7098 7935 7100
rect 7959 7098 8015 7100
rect 8039 7098 8095 7100
rect 8119 7098 8175 7100
rect 7879 7046 7925 7098
rect 7925 7046 7935 7098
rect 7959 7046 7989 7098
rect 7989 7046 8001 7098
rect 8001 7046 8015 7098
rect 8039 7046 8053 7098
rect 8053 7046 8065 7098
rect 8065 7046 8095 7098
rect 8119 7046 8129 7098
rect 8129 7046 8175 7098
rect 7879 7044 7935 7046
rect 7959 7044 8015 7046
rect 8039 7044 8095 7046
rect 8119 7044 8175 7046
rect 6561 6554 6617 6556
rect 6641 6554 6697 6556
rect 6721 6554 6777 6556
rect 6801 6554 6857 6556
rect 6561 6502 6607 6554
rect 6607 6502 6617 6554
rect 6641 6502 6671 6554
rect 6671 6502 6683 6554
rect 6683 6502 6697 6554
rect 6721 6502 6735 6554
rect 6735 6502 6747 6554
rect 6747 6502 6777 6554
rect 6801 6502 6811 6554
rect 6811 6502 6857 6554
rect 6561 6500 6617 6502
rect 6641 6500 6697 6502
rect 6721 6500 6777 6502
rect 6801 6500 6857 6502
rect 6550 5652 6552 5672
rect 6552 5652 6604 5672
rect 6604 5652 6606 5672
rect 6550 5616 6606 5652
rect 6561 5466 6617 5468
rect 6641 5466 6697 5468
rect 6721 5466 6777 5468
rect 6801 5466 6857 5468
rect 6561 5414 6607 5466
rect 6607 5414 6617 5466
rect 6641 5414 6671 5466
rect 6671 5414 6683 5466
rect 6683 5414 6697 5466
rect 6721 5414 6735 5466
rect 6735 5414 6747 5466
rect 6747 5414 6777 5466
rect 6801 5414 6811 5466
rect 6811 5414 6857 5466
rect 6561 5412 6617 5414
rect 6641 5412 6697 5414
rect 6721 5412 6777 5414
rect 6801 5412 6857 5414
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 4583 2202 4639 2204
rect 4663 2202 4719 2204
rect 4743 2202 4799 2204
rect 4823 2202 4879 2204
rect 4583 2150 4629 2202
rect 4629 2150 4639 2202
rect 4663 2150 4693 2202
rect 4693 2150 4705 2202
rect 4705 2150 4719 2202
rect 4743 2150 4757 2202
rect 4757 2150 4769 2202
rect 4769 2150 4799 2202
rect 4823 2150 4833 2202
rect 4833 2150 4879 2202
rect 4583 2148 4639 2150
rect 4663 2148 4719 2150
rect 4743 2148 4799 2150
rect 4823 2148 4879 2150
rect 5901 3834 5957 3836
rect 5981 3834 6037 3836
rect 6061 3834 6117 3836
rect 6141 3834 6197 3836
rect 5901 3782 5947 3834
rect 5947 3782 5957 3834
rect 5981 3782 6011 3834
rect 6011 3782 6023 3834
rect 6023 3782 6037 3834
rect 6061 3782 6075 3834
rect 6075 3782 6087 3834
rect 6087 3782 6117 3834
rect 6141 3782 6151 3834
rect 6151 3782 6197 3834
rect 5901 3780 5957 3782
rect 5981 3780 6037 3782
rect 6061 3780 6117 3782
rect 6141 3780 6197 3782
rect 5901 2746 5957 2748
rect 5981 2746 6037 2748
rect 6061 2746 6117 2748
rect 6141 2746 6197 2748
rect 5901 2694 5947 2746
rect 5947 2694 5957 2746
rect 5981 2694 6011 2746
rect 6011 2694 6023 2746
rect 6023 2694 6037 2746
rect 6061 2694 6075 2746
rect 6075 2694 6087 2746
rect 6087 2694 6117 2746
rect 6141 2694 6151 2746
rect 6151 2694 6197 2746
rect 5901 2692 5957 2694
rect 5981 2692 6037 2694
rect 6061 2692 6117 2694
rect 6141 2692 6197 2694
rect 6561 4378 6617 4380
rect 6641 4378 6697 4380
rect 6721 4378 6777 4380
rect 6801 4378 6857 4380
rect 6561 4326 6607 4378
rect 6607 4326 6617 4378
rect 6641 4326 6671 4378
rect 6671 4326 6683 4378
rect 6683 4326 6697 4378
rect 6721 4326 6735 4378
rect 6735 4326 6747 4378
rect 6747 4326 6777 4378
rect 6801 4326 6811 4378
rect 6811 4326 6857 4378
rect 6561 4324 6617 4326
rect 6641 4324 6697 4326
rect 6721 4324 6777 4326
rect 6801 4324 6857 4326
rect 7010 4120 7066 4176
rect 6561 3290 6617 3292
rect 6641 3290 6697 3292
rect 6721 3290 6777 3292
rect 6801 3290 6857 3292
rect 6561 3238 6607 3290
rect 6607 3238 6617 3290
rect 6641 3238 6671 3290
rect 6671 3238 6683 3290
rect 6683 3238 6697 3290
rect 6721 3238 6735 3290
rect 6735 3238 6747 3290
rect 6747 3238 6777 3290
rect 6801 3238 6811 3290
rect 6811 3238 6857 3290
rect 6561 3236 6617 3238
rect 6641 3236 6697 3238
rect 6721 3236 6777 3238
rect 6801 3236 6857 3238
rect 5998 1980 6000 2000
rect 6000 1980 6052 2000
rect 6052 1980 6054 2000
rect 5998 1944 6054 1980
rect 7879 6010 7935 6012
rect 7959 6010 8015 6012
rect 8039 6010 8095 6012
rect 8119 6010 8175 6012
rect 7879 5958 7925 6010
rect 7925 5958 7935 6010
rect 7959 5958 7989 6010
rect 7989 5958 8001 6010
rect 8001 5958 8015 6010
rect 8039 5958 8053 6010
rect 8053 5958 8065 6010
rect 8065 5958 8095 6010
rect 8119 5958 8129 6010
rect 8129 5958 8175 6010
rect 7879 5956 7935 5958
rect 7959 5956 8015 5958
rect 8039 5956 8095 5958
rect 8119 5956 8175 5958
rect 8539 8730 8595 8732
rect 8619 8730 8675 8732
rect 8699 8730 8755 8732
rect 8779 8730 8835 8732
rect 8539 8678 8585 8730
rect 8585 8678 8595 8730
rect 8619 8678 8649 8730
rect 8649 8678 8661 8730
rect 8661 8678 8675 8730
rect 8699 8678 8713 8730
rect 8713 8678 8725 8730
rect 8725 8678 8755 8730
rect 8779 8678 8789 8730
rect 8789 8678 8835 8730
rect 8539 8676 8595 8678
rect 8619 8676 8675 8678
rect 8699 8676 8755 8678
rect 8779 8676 8835 8678
rect 8942 8200 8998 8256
rect 8539 7642 8595 7644
rect 8619 7642 8675 7644
rect 8699 7642 8755 7644
rect 8779 7642 8835 7644
rect 8539 7590 8585 7642
rect 8585 7590 8595 7642
rect 8619 7590 8649 7642
rect 8649 7590 8661 7642
rect 8661 7590 8675 7642
rect 8699 7590 8713 7642
rect 8713 7590 8725 7642
rect 8725 7590 8755 7642
rect 8779 7590 8789 7642
rect 8789 7590 8835 7642
rect 8539 7588 8595 7590
rect 8619 7588 8675 7590
rect 8699 7588 8755 7590
rect 8779 7588 8835 7590
rect 8942 7520 8998 7576
rect 7879 4922 7935 4924
rect 7959 4922 8015 4924
rect 8039 4922 8095 4924
rect 8119 4922 8175 4924
rect 7879 4870 7925 4922
rect 7925 4870 7935 4922
rect 7959 4870 7989 4922
rect 7989 4870 8001 4922
rect 8001 4870 8015 4922
rect 8039 4870 8053 4922
rect 8053 4870 8065 4922
rect 8065 4870 8095 4922
rect 8119 4870 8129 4922
rect 8129 4870 8175 4922
rect 7879 4868 7935 4870
rect 7959 4868 8015 4870
rect 8039 4868 8095 4870
rect 8119 4868 8175 4870
rect 8574 6840 8630 6896
rect 8539 6554 8595 6556
rect 8619 6554 8675 6556
rect 8699 6554 8755 6556
rect 8779 6554 8835 6556
rect 8539 6502 8585 6554
rect 8585 6502 8595 6554
rect 8619 6502 8649 6554
rect 8649 6502 8661 6554
rect 8661 6502 8675 6554
rect 8699 6502 8713 6554
rect 8713 6502 8725 6554
rect 8725 6502 8755 6554
rect 8779 6502 8789 6554
rect 8789 6502 8835 6554
rect 8539 6500 8595 6502
rect 8619 6500 8675 6502
rect 8699 6500 8755 6502
rect 8779 6500 8835 6502
rect 8574 6160 8630 6216
rect 9126 7384 9182 7440
rect 8942 5480 8998 5536
rect 8539 5466 8595 5468
rect 8619 5466 8675 5468
rect 8699 5466 8755 5468
rect 8779 5466 8835 5468
rect 8539 5414 8585 5466
rect 8585 5414 8595 5466
rect 8619 5414 8649 5466
rect 8649 5414 8661 5466
rect 8661 5414 8675 5466
rect 8699 5414 8713 5466
rect 8713 5414 8725 5466
rect 8725 5414 8755 5466
rect 8779 5414 8789 5466
rect 8789 5414 8835 5466
rect 8539 5412 8595 5414
rect 8619 5412 8675 5414
rect 8699 5412 8755 5414
rect 8779 5412 8835 5414
rect 8539 4378 8595 4380
rect 8619 4378 8675 4380
rect 8699 4378 8755 4380
rect 8779 4378 8835 4380
rect 8539 4326 8585 4378
rect 8585 4326 8595 4378
rect 8619 4326 8649 4378
rect 8649 4326 8661 4378
rect 8661 4326 8675 4378
rect 8699 4326 8713 4378
rect 8713 4326 8725 4378
rect 8725 4326 8755 4378
rect 8779 4326 8789 4378
rect 8789 4326 8835 4378
rect 8539 4324 8595 4326
rect 8619 4324 8675 4326
rect 8699 4324 8755 4326
rect 8779 4324 8835 4326
rect 7879 3834 7935 3836
rect 7959 3834 8015 3836
rect 8039 3834 8095 3836
rect 8119 3834 8175 3836
rect 7879 3782 7925 3834
rect 7925 3782 7935 3834
rect 7959 3782 7989 3834
rect 7989 3782 8001 3834
rect 8001 3782 8015 3834
rect 8039 3782 8053 3834
rect 8053 3782 8065 3834
rect 8065 3782 8095 3834
rect 8119 3782 8129 3834
rect 8129 3782 8175 3834
rect 7879 3780 7935 3782
rect 7959 3780 8015 3782
rect 8039 3780 8095 3782
rect 8119 3780 8175 3782
rect 7378 2760 7434 2816
rect 8482 3440 8538 3496
rect 7746 2760 7802 2816
rect 7879 2746 7935 2748
rect 7959 2746 8015 2748
rect 8039 2746 8095 2748
rect 8119 2746 8175 2748
rect 7879 2694 7925 2746
rect 7925 2694 7935 2746
rect 7959 2694 7989 2746
rect 7989 2694 8001 2746
rect 8001 2694 8015 2746
rect 8039 2694 8053 2746
rect 8053 2694 8065 2746
rect 8065 2694 8095 2746
rect 8119 2694 8129 2746
rect 8129 2694 8175 2746
rect 7879 2692 7935 2694
rect 7959 2692 8015 2694
rect 8039 2692 8095 2694
rect 8119 2692 8175 2694
rect 8539 3290 8595 3292
rect 8619 3290 8675 3292
rect 8699 3290 8755 3292
rect 8779 3290 8835 3292
rect 8539 3238 8585 3290
rect 8585 3238 8595 3290
rect 8619 3238 8649 3290
rect 8649 3238 8661 3290
rect 8661 3238 8675 3290
rect 8699 3238 8713 3290
rect 8713 3238 8725 3290
rect 8725 3238 8755 3290
rect 8779 3238 8789 3290
rect 8789 3238 8835 3290
rect 8539 3236 8595 3238
rect 8619 3236 8675 3238
rect 8699 3236 8755 3238
rect 8779 3236 8835 3238
rect 6561 2202 6617 2204
rect 6641 2202 6697 2204
rect 6721 2202 6777 2204
rect 6801 2202 6857 2204
rect 6561 2150 6607 2202
rect 6607 2150 6617 2202
rect 6641 2150 6671 2202
rect 6671 2150 6683 2202
rect 6683 2150 6697 2202
rect 6721 2150 6735 2202
rect 6735 2150 6747 2202
rect 6747 2150 6777 2202
rect 6801 2150 6811 2202
rect 6811 2150 6857 2202
rect 6561 2148 6617 2150
rect 6641 2148 6697 2150
rect 6721 2148 6777 2150
rect 6801 2148 6857 2150
rect 8539 2202 8595 2204
rect 8619 2202 8675 2204
rect 8699 2202 8755 2204
rect 8779 2202 8835 2204
rect 8539 2150 8585 2202
rect 8585 2150 8595 2202
rect 8619 2150 8649 2202
rect 8649 2150 8661 2202
rect 8661 2150 8675 2202
rect 8699 2150 8713 2202
rect 8713 2150 8725 2202
rect 8725 2150 8755 2202
rect 8779 2150 8789 2202
rect 8789 2150 8835 2202
rect 8539 2148 8595 2150
rect 8619 2148 8675 2150
rect 8699 2148 8755 2150
rect 8779 2148 8835 2150
<< metal3 >>
rect 2595 9824 2911 9825
rect 2595 9760 2601 9824
rect 2665 9760 2681 9824
rect 2745 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2911 9824
rect 2595 9759 2911 9760
rect 4573 9824 4889 9825
rect 4573 9760 4579 9824
rect 4643 9760 4659 9824
rect 4723 9760 4739 9824
rect 4803 9760 4819 9824
rect 4883 9760 4889 9824
rect 4573 9759 4889 9760
rect 6551 9824 6867 9825
rect 6551 9760 6557 9824
rect 6621 9760 6637 9824
rect 6701 9760 6717 9824
rect 6781 9760 6797 9824
rect 6861 9760 6867 9824
rect 6551 9759 6867 9760
rect 8529 9824 8845 9825
rect 8529 9760 8535 9824
rect 8599 9760 8615 9824
rect 8679 9760 8695 9824
rect 8759 9760 8775 9824
rect 8839 9760 8845 9824
rect 8529 9759 8845 9760
rect 0 9618 800 9648
rect 1025 9618 1091 9621
rect 0 9616 1091 9618
rect 0 9560 1030 9616
rect 1086 9560 1091 9616
rect 0 9558 1091 9560
rect 0 9528 800 9558
rect 1025 9555 1091 9558
rect 1935 9280 2251 9281
rect 1935 9216 1941 9280
rect 2005 9216 2021 9280
rect 2085 9216 2101 9280
rect 2165 9216 2181 9280
rect 2245 9216 2251 9280
rect 1935 9215 2251 9216
rect 3913 9280 4229 9281
rect 3913 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4229 9280
rect 3913 9215 4229 9216
rect 5891 9280 6207 9281
rect 5891 9216 5897 9280
rect 5961 9216 5977 9280
rect 6041 9216 6057 9280
rect 6121 9216 6137 9280
rect 6201 9216 6207 9280
rect 5891 9215 6207 9216
rect 7869 9280 8185 9281
rect 7869 9216 7875 9280
rect 7939 9216 7955 9280
rect 8019 9216 8035 9280
rect 8099 9216 8115 9280
rect 8179 9216 8185 9280
rect 7869 9215 8185 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 7005 8938 7071 8941
rect 9401 8938 10201 8968
rect 7005 8936 10201 8938
rect 7005 8880 7010 8936
rect 7066 8880 10201 8936
rect 7005 8878 10201 8880
rect 7005 8875 7071 8878
rect 9401 8848 10201 8878
rect 2595 8736 2911 8737
rect 2595 8672 2601 8736
rect 2665 8672 2681 8736
rect 2745 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2911 8736
rect 2595 8671 2911 8672
rect 4573 8736 4889 8737
rect 4573 8672 4579 8736
rect 4643 8672 4659 8736
rect 4723 8672 4739 8736
rect 4803 8672 4819 8736
rect 4883 8672 4889 8736
rect 4573 8671 4889 8672
rect 6551 8736 6867 8737
rect 6551 8672 6557 8736
rect 6621 8672 6637 8736
rect 6701 8672 6717 8736
rect 6781 8672 6797 8736
rect 6861 8672 6867 8736
rect 6551 8671 6867 8672
rect 8529 8736 8845 8737
rect 8529 8672 8535 8736
rect 8599 8672 8615 8736
rect 8679 8672 8695 8736
rect 8759 8672 8775 8736
rect 8839 8672 8845 8736
rect 8529 8671 8845 8672
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 8937 8258 9003 8261
rect 9401 8258 10201 8288
rect 8937 8256 10201 8258
rect 8937 8200 8942 8256
rect 8998 8200 10201 8256
rect 8937 8198 10201 8200
rect 8937 8195 9003 8198
rect 1935 8192 2251 8193
rect 1935 8128 1941 8192
rect 2005 8128 2021 8192
rect 2085 8128 2101 8192
rect 2165 8128 2181 8192
rect 2245 8128 2251 8192
rect 1935 8127 2251 8128
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 5891 8192 6207 8193
rect 5891 8128 5897 8192
rect 5961 8128 5977 8192
rect 6041 8128 6057 8192
rect 6121 8128 6137 8192
rect 6201 8128 6207 8192
rect 5891 8127 6207 8128
rect 7869 8192 8185 8193
rect 7869 8128 7875 8192
rect 7939 8128 7955 8192
rect 8019 8128 8035 8192
rect 8099 8128 8115 8192
rect 8179 8128 8185 8192
rect 9401 8168 10201 8198
rect 7869 8127 8185 8128
rect 2595 7648 2911 7649
rect 0 7578 800 7608
rect 2595 7584 2601 7648
rect 2665 7584 2681 7648
rect 2745 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2911 7648
rect 2595 7583 2911 7584
rect 4573 7648 4889 7649
rect 4573 7584 4579 7648
rect 4643 7584 4659 7648
rect 4723 7584 4739 7648
rect 4803 7584 4819 7648
rect 4883 7584 4889 7648
rect 4573 7583 4889 7584
rect 6551 7648 6867 7649
rect 6551 7584 6557 7648
rect 6621 7584 6637 7648
rect 6701 7584 6717 7648
rect 6781 7584 6797 7648
rect 6861 7584 6867 7648
rect 6551 7583 6867 7584
rect 8529 7648 8845 7649
rect 8529 7584 8535 7648
rect 8599 7584 8615 7648
rect 8679 7584 8695 7648
rect 8759 7584 8775 7648
rect 8839 7584 8845 7648
rect 8529 7583 8845 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 8937 7578 9003 7581
rect 9401 7578 10201 7608
rect 8937 7576 10201 7578
rect 8937 7520 8942 7576
rect 8998 7520 10201 7576
rect 8937 7518 10201 7520
rect 8937 7515 9003 7518
rect 9401 7488 10201 7518
rect 6729 7442 6795 7445
rect 9121 7442 9187 7445
rect 6729 7440 9187 7442
rect 6729 7384 6734 7440
rect 6790 7384 9126 7440
rect 9182 7384 9187 7440
rect 6729 7382 9187 7384
rect 6729 7379 6795 7382
rect 9121 7379 9187 7382
rect 5349 7306 5415 7309
rect 7557 7306 7623 7309
rect 5349 7304 7623 7306
rect 5349 7248 5354 7304
rect 5410 7248 7562 7304
rect 7618 7248 7623 7304
rect 5349 7246 7623 7248
rect 5349 7243 5415 7246
rect 7557 7243 7623 7246
rect 1935 7104 2251 7105
rect 1935 7040 1941 7104
rect 2005 7040 2021 7104
rect 2085 7040 2101 7104
rect 2165 7040 2181 7104
rect 2245 7040 2251 7104
rect 1935 7039 2251 7040
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 5891 7104 6207 7105
rect 5891 7040 5897 7104
rect 5961 7040 5977 7104
rect 6041 7040 6057 7104
rect 6121 7040 6137 7104
rect 6201 7040 6207 7104
rect 5891 7039 6207 7040
rect 7869 7104 8185 7105
rect 7869 7040 7875 7104
rect 7939 7040 7955 7104
rect 8019 7040 8035 7104
rect 8099 7040 8115 7104
rect 8179 7040 8185 7104
rect 7869 7039 8185 7040
rect 0 6900 800 6928
rect 0 6836 796 6900
rect 860 6836 866 6900
rect 8569 6898 8635 6901
rect 9401 6898 10201 6928
rect 8569 6896 10201 6898
rect 8569 6840 8574 6896
rect 8630 6840 10201 6896
rect 8569 6838 10201 6840
rect 0 6808 800 6836
rect 8569 6835 8635 6838
rect 9401 6808 10201 6838
rect 841 6628 907 6629
rect 790 6626 796 6628
rect 750 6566 796 6626
rect 860 6624 907 6628
rect 902 6568 907 6624
rect 790 6564 796 6566
rect 860 6564 907 6568
rect 841 6563 907 6564
rect 2595 6560 2911 6561
rect 2595 6496 2601 6560
rect 2665 6496 2681 6560
rect 2745 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2911 6560
rect 2595 6495 2911 6496
rect 4573 6560 4889 6561
rect 4573 6496 4579 6560
rect 4643 6496 4659 6560
rect 4723 6496 4739 6560
rect 4803 6496 4819 6560
rect 4883 6496 4889 6560
rect 4573 6495 4889 6496
rect 6551 6560 6867 6561
rect 6551 6496 6557 6560
rect 6621 6496 6637 6560
rect 6701 6496 6717 6560
rect 6781 6496 6797 6560
rect 6861 6496 6867 6560
rect 6551 6495 6867 6496
rect 8529 6560 8845 6561
rect 8529 6496 8535 6560
rect 8599 6496 8615 6560
rect 8679 6496 8695 6560
rect 8759 6496 8775 6560
rect 8839 6496 8845 6560
rect 8529 6495 8845 6496
rect 0 6220 800 6248
rect 0 6156 796 6220
rect 860 6156 866 6220
rect 8569 6218 8635 6221
rect 9401 6218 10201 6248
rect 8569 6216 10201 6218
rect 8569 6160 8574 6216
rect 8630 6160 10201 6216
rect 8569 6158 10201 6160
rect 0 6128 800 6156
rect 8569 6155 8635 6158
rect 9401 6128 10201 6158
rect 1935 6016 2251 6017
rect 1935 5952 1941 6016
rect 2005 5952 2021 6016
rect 2085 5952 2101 6016
rect 2165 5952 2181 6016
rect 2245 5952 2251 6016
rect 1935 5951 2251 5952
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 5891 6016 6207 6017
rect 5891 5952 5897 6016
rect 5961 5952 5977 6016
rect 6041 5952 6057 6016
rect 6121 5952 6137 6016
rect 6201 5952 6207 6016
rect 5891 5951 6207 5952
rect 7869 6016 8185 6017
rect 7869 5952 7875 6016
rect 7939 5952 7955 6016
rect 8019 5952 8035 6016
rect 8099 5952 8115 6016
rect 8179 5952 8185 6016
rect 7869 5951 8185 5952
rect 841 5948 907 5949
rect 790 5946 796 5948
rect 750 5886 796 5946
rect 860 5944 907 5948
rect 902 5888 907 5944
rect 790 5884 796 5886
rect 860 5884 907 5888
rect 841 5883 907 5884
rect 1393 5810 1459 5813
rect 4337 5810 4403 5813
rect 1393 5808 4403 5810
rect 1393 5752 1398 5808
rect 1454 5752 4342 5808
rect 4398 5752 4403 5808
rect 1393 5750 4403 5752
rect 1393 5747 1459 5750
rect 4337 5747 4403 5750
rect 5073 5674 5139 5677
rect 6545 5674 6611 5677
rect 5073 5672 6611 5674
rect 5073 5616 5078 5672
rect 5134 5616 6550 5672
rect 6606 5616 6611 5672
rect 5073 5614 6611 5616
rect 5073 5611 5139 5614
rect 6545 5611 6611 5614
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 8937 5538 9003 5541
rect 9401 5538 10201 5568
rect 8937 5536 10201 5538
rect 8937 5480 8942 5536
rect 8998 5480 10201 5536
rect 8937 5478 10201 5480
rect 8937 5475 9003 5478
rect 2595 5472 2911 5473
rect 2595 5408 2601 5472
rect 2665 5408 2681 5472
rect 2745 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2911 5472
rect 2595 5407 2911 5408
rect 4573 5472 4889 5473
rect 4573 5408 4579 5472
rect 4643 5408 4659 5472
rect 4723 5408 4739 5472
rect 4803 5408 4819 5472
rect 4883 5408 4889 5472
rect 4573 5407 4889 5408
rect 6551 5472 6867 5473
rect 6551 5408 6557 5472
rect 6621 5408 6637 5472
rect 6701 5408 6717 5472
rect 6781 5408 6797 5472
rect 6861 5408 6867 5472
rect 6551 5407 6867 5408
rect 8529 5472 8845 5473
rect 8529 5408 8535 5472
rect 8599 5408 8615 5472
rect 8679 5408 8695 5472
rect 8759 5408 8775 5472
rect 8839 5408 8845 5472
rect 9401 5448 10201 5478
rect 8529 5407 8845 5408
rect 5717 5266 5783 5269
rect 6085 5266 6151 5269
rect 5717 5264 6151 5266
rect 5717 5208 5722 5264
rect 5778 5208 6090 5264
rect 6146 5208 6151 5264
rect 5717 5206 6151 5208
rect 5717 5203 5783 5206
rect 6085 5203 6151 5206
rect 5349 4994 5415 4997
rect 5349 4992 5458 4994
rect 5349 4936 5354 4992
rect 5410 4936 5458 4992
rect 5349 4931 5458 4936
rect 1935 4928 2251 4929
rect 0 4858 800 4888
rect 1935 4864 1941 4928
rect 2005 4864 2021 4928
rect 2085 4864 2101 4928
rect 2165 4864 2181 4928
rect 2245 4864 2251 4928
rect 1935 4863 2251 4864
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 5398 4725 5458 4931
rect 5891 4928 6207 4929
rect 5891 4864 5897 4928
rect 5961 4864 5977 4928
rect 6041 4864 6057 4928
rect 6121 4864 6137 4928
rect 6201 4864 6207 4928
rect 5891 4863 6207 4864
rect 7869 4928 8185 4929
rect 7869 4864 7875 4928
rect 7939 4864 7955 4928
rect 8019 4864 8035 4928
rect 8099 4864 8115 4928
rect 8179 4864 8185 4928
rect 7869 4863 8185 4864
rect 9401 4858 10201 4888
rect 8342 4798 10201 4858
rect 5349 4720 5458 4725
rect 5349 4664 5354 4720
rect 5410 4664 5458 4720
rect 5349 4662 5458 4664
rect 6177 4722 6243 4725
rect 8342 4722 8402 4798
rect 9401 4768 10201 4798
rect 6177 4720 8402 4722
rect 6177 4664 6182 4720
rect 6238 4664 8402 4720
rect 6177 4662 8402 4664
rect 5349 4659 5415 4662
rect 6177 4659 6243 4662
rect 2595 4384 2911 4385
rect 2595 4320 2601 4384
rect 2665 4320 2681 4384
rect 2745 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2911 4384
rect 2595 4319 2911 4320
rect 4573 4384 4889 4385
rect 4573 4320 4579 4384
rect 4643 4320 4659 4384
rect 4723 4320 4739 4384
rect 4803 4320 4819 4384
rect 4883 4320 4889 4384
rect 4573 4319 4889 4320
rect 6551 4384 6867 4385
rect 6551 4320 6557 4384
rect 6621 4320 6637 4384
rect 6701 4320 6717 4384
rect 6781 4320 6797 4384
rect 6861 4320 6867 4384
rect 6551 4319 6867 4320
rect 8529 4384 8845 4385
rect 8529 4320 8535 4384
rect 8599 4320 8615 4384
rect 8679 4320 8695 4384
rect 8759 4320 8775 4384
rect 8839 4320 8845 4384
rect 8529 4319 8845 4320
rect 7005 4178 7071 4181
rect 9401 4178 10201 4208
rect 7005 4176 10201 4178
rect 7005 4120 7010 4176
rect 7066 4120 10201 4176
rect 7005 4118 10201 4120
rect 7005 4115 7071 4118
rect 9401 4088 10201 4118
rect 1935 3840 2251 3841
rect 1935 3776 1941 3840
rect 2005 3776 2021 3840
rect 2085 3776 2101 3840
rect 2165 3776 2181 3840
rect 2245 3776 2251 3840
rect 1935 3775 2251 3776
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 5891 3840 6207 3841
rect 5891 3776 5897 3840
rect 5961 3776 5977 3840
rect 6041 3776 6057 3840
rect 6121 3776 6137 3840
rect 6201 3776 6207 3840
rect 5891 3775 6207 3776
rect 7869 3840 8185 3841
rect 7869 3776 7875 3840
rect 7939 3776 7955 3840
rect 8019 3776 8035 3840
rect 8099 3776 8115 3840
rect 8179 3776 8185 3840
rect 7869 3775 8185 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 8477 3498 8543 3501
rect 9401 3498 10201 3528
rect 8477 3496 10201 3498
rect 8477 3440 8482 3496
rect 8538 3440 10201 3496
rect 8477 3438 10201 3440
rect 8477 3435 8543 3438
rect 9401 3408 10201 3438
rect 2595 3296 2911 3297
rect 2595 3232 2601 3296
rect 2665 3232 2681 3296
rect 2745 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2911 3296
rect 2595 3231 2911 3232
rect 4573 3296 4889 3297
rect 4573 3232 4579 3296
rect 4643 3232 4659 3296
rect 4723 3232 4739 3296
rect 4803 3232 4819 3296
rect 4883 3232 4889 3296
rect 4573 3231 4889 3232
rect 6551 3296 6867 3297
rect 6551 3232 6557 3296
rect 6621 3232 6637 3296
rect 6701 3232 6717 3296
rect 6781 3232 6797 3296
rect 6861 3232 6867 3296
rect 6551 3231 6867 3232
rect 8529 3296 8845 3297
rect 8529 3232 8535 3296
rect 8599 3232 8615 3296
rect 8679 3232 8695 3296
rect 8759 3232 8775 3296
rect 8839 3232 8845 3296
rect 8529 3231 8845 3232
rect 7373 2818 7439 2821
rect 7741 2818 7807 2821
rect 9401 2818 10201 2848
rect 7373 2816 7807 2818
rect 7373 2760 7378 2816
rect 7434 2760 7746 2816
rect 7802 2760 7807 2816
rect 7373 2758 7807 2760
rect 7373 2755 7439 2758
rect 7741 2755 7807 2758
rect 8342 2758 10201 2818
rect 1935 2752 2251 2753
rect 1935 2688 1941 2752
rect 2005 2688 2021 2752
rect 2085 2688 2101 2752
rect 2165 2688 2181 2752
rect 2245 2688 2251 2752
rect 1935 2687 2251 2688
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 5891 2752 6207 2753
rect 5891 2688 5897 2752
rect 5961 2688 5977 2752
rect 6041 2688 6057 2752
rect 6121 2688 6137 2752
rect 6201 2688 6207 2752
rect 5891 2687 6207 2688
rect 7869 2752 8185 2753
rect 7869 2688 7875 2752
rect 7939 2688 7955 2752
rect 8019 2688 8035 2752
rect 8099 2688 8115 2752
rect 8179 2688 8185 2752
rect 7869 2687 8185 2688
rect 1669 2546 1735 2549
rect 8342 2546 8402 2758
rect 9401 2728 10201 2758
rect 1669 2544 8402 2546
rect 1669 2488 1674 2544
rect 1730 2488 8402 2544
rect 1669 2486 8402 2488
rect 1669 2483 1735 2486
rect 2595 2208 2911 2209
rect 2595 2144 2601 2208
rect 2665 2144 2681 2208
rect 2745 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2911 2208
rect 2595 2143 2911 2144
rect 4573 2208 4889 2209
rect 4573 2144 4579 2208
rect 4643 2144 4659 2208
rect 4723 2144 4739 2208
rect 4803 2144 4819 2208
rect 4883 2144 4889 2208
rect 4573 2143 4889 2144
rect 6551 2208 6867 2209
rect 6551 2144 6557 2208
rect 6621 2144 6637 2208
rect 6701 2144 6717 2208
rect 6781 2144 6797 2208
rect 6861 2144 6867 2208
rect 6551 2143 6867 2144
rect 8529 2208 8845 2209
rect 8529 2144 8535 2208
rect 8599 2144 8615 2208
rect 8679 2144 8695 2208
rect 8759 2144 8775 2208
rect 8839 2144 8845 2208
rect 8529 2143 8845 2144
rect 9401 2138 10201 2168
rect 9078 2078 10201 2138
rect 5993 2002 6059 2005
rect 9078 2002 9138 2078
rect 9401 2048 10201 2078
rect 5993 2000 9138 2002
rect 5993 1944 5998 2000
rect 6054 1944 9138 2000
rect 5993 1942 9138 1944
rect 5993 1939 6059 1942
<< via3 >>
rect 2601 9820 2665 9824
rect 2601 9764 2605 9820
rect 2605 9764 2661 9820
rect 2661 9764 2665 9820
rect 2601 9760 2665 9764
rect 2681 9820 2745 9824
rect 2681 9764 2685 9820
rect 2685 9764 2741 9820
rect 2741 9764 2745 9820
rect 2681 9760 2745 9764
rect 2761 9820 2825 9824
rect 2761 9764 2765 9820
rect 2765 9764 2821 9820
rect 2821 9764 2825 9820
rect 2761 9760 2825 9764
rect 2841 9820 2905 9824
rect 2841 9764 2845 9820
rect 2845 9764 2901 9820
rect 2901 9764 2905 9820
rect 2841 9760 2905 9764
rect 4579 9820 4643 9824
rect 4579 9764 4583 9820
rect 4583 9764 4639 9820
rect 4639 9764 4643 9820
rect 4579 9760 4643 9764
rect 4659 9820 4723 9824
rect 4659 9764 4663 9820
rect 4663 9764 4719 9820
rect 4719 9764 4723 9820
rect 4659 9760 4723 9764
rect 4739 9820 4803 9824
rect 4739 9764 4743 9820
rect 4743 9764 4799 9820
rect 4799 9764 4803 9820
rect 4739 9760 4803 9764
rect 4819 9820 4883 9824
rect 4819 9764 4823 9820
rect 4823 9764 4879 9820
rect 4879 9764 4883 9820
rect 4819 9760 4883 9764
rect 6557 9820 6621 9824
rect 6557 9764 6561 9820
rect 6561 9764 6617 9820
rect 6617 9764 6621 9820
rect 6557 9760 6621 9764
rect 6637 9820 6701 9824
rect 6637 9764 6641 9820
rect 6641 9764 6697 9820
rect 6697 9764 6701 9820
rect 6637 9760 6701 9764
rect 6717 9820 6781 9824
rect 6717 9764 6721 9820
rect 6721 9764 6777 9820
rect 6777 9764 6781 9820
rect 6717 9760 6781 9764
rect 6797 9820 6861 9824
rect 6797 9764 6801 9820
rect 6801 9764 6857 9820
rect 6857 9764 6861 9820
rect 6797 9760 6861 9764
rect 8535 9820 8599 9824
rect 8535 9764 8539 9820
rect 8539 9764 8595 9820
rect 8595 9764 8599 9820
rect 8535 9760 8599 9764
rect 8615 9820 8679 9824
rect 8615 9764 8619 9820
rect 8619 9764 8675 9820
rect 8675 9764 8679 9820
rect 8615 9760 8679 9764
rect 8695 9820 8759 9824
rect 8695 9764 8699 9820
rect 8699 9764 8755 9820
rect 8755 9764 8759 9820
rect 8695 9760 8759 9764
rect 8775 9820 8839 9824
rect 8775 9764 8779 9820
rect 8779 9764 8835 9820
rect 8835 9764 8839 9820
rect 8775 9760 8839 9764
rect 1941 9276 2005 9280
rect 1941 9220 1945 9276
rect 1945 9220 2001 9276
rect 2001 9220 2005 9276
rect 1941 9216 2005 9220
rect 2021 9276 2085 9280
rect 2021 9220 2025 9276
rect 2025 9220 2081 9276
rect 2081 9220 2085 9276
rect 2021 9216 2085 9220
rect 2101 9276 2165 9280
rect 2101 9220 2105 9276
rect 2105 9220 2161 9276
rect 2161 9220 2165 9276
rect 2101 9216 2165 9220
rect 2181 9276 2245 9280
rect 2181 9220 2185 9276
rect 2185 9220 2241 9276
rect 2241 9220 2245 9276
rect 2181 9216 2245 9220
rect 3919 9276 3983 9280
rect 3919 9220 3923 9276
rect 3923 9220 3979 9276
rect 3979 9220 3983 9276
rect 3919 9216 3983 9220
rect 3999 9276 4063 9280
rect 3999 9220 4003 9276
rect 4003 9220 4059 9276
rect 4059 9220 4063 9276
rect 3999 9216 4063 9220
rect 4079 9276 4143 9280
rect 4079 9220 4083 9276
rect 4083 9220 4139 9276
rect 4139 9220 4143 9276
rect 4079 9216 4143 9220
rect 4159 9276 4223 9280
rect 4159 9220 4163 9276
rect 4163 9220 4219 9276
rect 4219 9220 4223 9276
rect 4159 9216 4223 9220
rect 5897 9276 5961 9280
rect 5897 9220 5901 9276
rect 5901 9220 5957 9276
rect 5957 9220 5961 9276
rect 5897 9216 5961 9220
rect 5977 9276 6041 9280
rect 5977 9220 5981 9276
rect 5981 9220 6037 9276
rect 6037 9220 6041 9276
rect 5977 9216 6041 9220
rect 6057 9276 6121 9280
rect 6057 9220 6061 9276
rect 6061 9220 6117 9276
rect 6117 9220 6121 9276
rect 6057 9216 6121 9220
rect 6137 9276 6201 9280
rect 6137 9220 6141 9276
rect 6141 9220 6197 9276
rect 6197 9220 6201 9276
rect 6137 9216 6201 9220
rect 7875 9276 7939 9280
rect 7875 9220 7879 9276
rect 7879 9220 7935 9276
rect 7935 9220 7939 9276
rect 7875 9216 7939 9220
rect 7955 9276 8019 9280
rect 7955 9220 7959 9276
rect 7959 9220 8015 9276
rect 8015 9220 8019 9276
rect 7955 9216 8019 9220
rect 8035 9276 8099 9280
rect 8035 9220 8039 9276
rect 8039 9220 8095 9276
rect 8095 9220 8099 9276
rect 8035 9216 8099 9220
rect 8115 9276 8179 9280
rect 8115 9220 8119 9276
rect 8119 9220 8175 9276
rect 8175 9220 8179 9276
rect 8115 9216 8179 9220
rect 2601 8732 2665 8736
rect 2601 8676 2605 8732
rect 2605 8676 2661 8732
rect 2661 8676 2665 8732
rect 2601 8672 2665 8676
rect 2681 8732 2745 8736
rect 2681 8676 2685 8732
rect 2685 8676 2741 8732
rect 2741 8676 2745 8732
rect 2681 8672 2745 8676
rect 2761 8732 2825 8736
rect 2761 8676 2765 8732
rect 2765 8676 2821 8732
rect 2821 8676 2825 8732
rect 2761 8672 2825 8676
rect 2841 8732 2905 8736
rect 2841 8676 2845 8732
rect 2845 8676 2901 8732
rect 2901 8676 2905 8732
rect 2841 8672 2905 8676
rect 4579 8732 4643 8736
rect 4579 8676 4583 8732
rect 4583 8676 4639 8732
rect 4639 8676 4643 8732
rect 4579 8672 4643 8676
rect 4659 8732 4723 8736
rect 4659 8676 4663 8732
rect 4663 8676 4719 8732
rect 4719 8676 4723 8732
rect 4659 8672 4723 8676
rect 4739 8732 4803 8736
rect 4739 8676 4743 8732
rect 4743 8676 4799 8732
rect 4799 8676 4803 8732
rect 4739 8672 4803 8676
rect 4819 8732 4883 8736
rect 4819 8676 4823 8732
rect 4823 8676 4879 8732
rect 4879 8676 4883 8732
rect 4819 8672 4883 8676
rect 6557 8732 6621 8736
rect 6557 8676 6561 8732
rect 6561 8676 6617 8732
rect 6617 8676 6621 8732
rect 6557 8672 6621 8676
rect 6637 8732 6701 8736
rect 6637 8676 6641 8732
rect 6641 8676 6697 8732
rect 6697 8676 6701 8732
rect 6637 8672 6701 8676
rect 6717 8732 6781 8736
rect 6717 8676 6721 8732
rect 6721 8676 6777 8732
rect 6777 8676 6781 8732
rect 6717 8672 6781 8676
rect 6797 8732 6861 8736
rect 6797 8676 6801 8732
rect 6801 8676 6857 8732
rect 6857 8676 6861 8732
rect 6797 8672 6861 8676
rect 8535 8732 8599 8736
rect 8535 8676 8539 8732
rect 8539 8676 8595 8732
rect 8595 8676 8599 8732
rect 8535 8672 8599 8676
rect 8615 8732 8679 8736
rect 8615 8676 8619 8732
rect 8619 8676 8675 8732
rect 8675 8676 8679 8732
rect 8615 8672 8679 8676
rect 8695 8732 8759 8736
rect 8695 8676 8699 8732
rect 8699 8676 8755 8732
rect 8755 8676 8759 8732
rect 8695 8672 8759 8676
rect 8775 8732 8839 8736
rect 8775 8676 8779 8732
rect 8779 8676 8835 8732
rect 8835 8676 8839 8732
rect 8775 8672 8839 8676
rect 1941 8188 2005 8192
rect 1941 8132 1945 8188
rect 1945 8132 2001 8188
rect 2001 8132 2005 8188
rect 1941 8128 2005 8132
rect 2021 8188 2085 8192
rect 2021 8132 2025 8188
rect 2025 8132 2081 8188
rect 2081 8132 2085 8188
rect 2021 8128 2085 8132
rect 2101 8188 2165 8192
rect 2101 8132 2105 8188
rect 2105 8132 2161 8188
rect 2161 8132 2165 8188
rect 2101 8128 2165 8132
rect 2181 8188 2245 8192
rect 2181 8132 2185 8188
rect 2185 8132 2241 8188
rect 2241 8132 2245 8188
rect 2181 8128 2245 8132
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 5897 8188 5961 8192
rect 5897 8132 5901 8188
rect 5901 8132 5957 8188
rect 5957 8132 5961 8188
rect 5897 8128 5961 8132
rect 5977 8188 6041 8192
rect 5977 8132 5981 8188
rect 5981 8132 6037 8188
rect 6037 8132 6041 8188
rect 5977 8128 6041 8132
rect 6057 8188 6121 8192
rect 6057 8132 6061 8188
rect 6061 8132 6117 8188
rect 6117 8132 6121 8188
rect 6057 8128 6121 8132
rect 6137 8188 6201 8192
rect 6137 8132 6141 8188
rect 6141 8132 6197 8188
rect 6197 8132 6201 8188
rect 6137 8128 6201 8132
rect 7875 8188 7939 8192
rect 7875 8132 7879 8188
rect 7879 8132 7935 8188
rect 7935 8132 7939 8188
rect 7875 8128 7939 8132
rect 7955 8188 8019 8192
rect 7955 8132 7959 8188
rect 7959 8132 8015 8188
rect 8015 8132 8019 8188
rect 7955 8128 8019 8132
rect 8035 8188 8099 8192
rect 8035 8132 8039 8188
rect 8039 8132 8095 8188
rect 8095 8132 8099 8188
rect 8035 8128 8099 8132
rect 8115 8188 8179 8192
rect 8115 8132 8119 8188
rect 8119 8132 8175 8188
rect 8175 8132 8179 8188
rect 8115 8128 8179 8132
rect 2601 7644 2665 7648
rect 2601 7588 2605 7644
rect 2605 7588 2661 7644
rect 2661 7588 2665 7644
rect 2601 7584 2665 7588
rect 2681 7644 2745 7648
rect 2681 7588 2685 7644
rect 2685 7588 2741 7644
rect 2741 7588 2745 7644
rect 2681 7584 2745 7588
rect 2761 7644 2825 7648
rect 2761 7588 2765 7644
rect 2765 7588 2821 7644
rect 2821 7588 2825 7644
rect 2761 7584 2825 7588
rect 2841 7644 2905 7648
rect 2841 7588 2845 7644
rect 2845 7588 2901 7644
rect 2901 7588 2905 7644
rect 2841 7584 2905 7588
rect 4579 7644 4643 7648
rect 4579 7588 4583 7644
rect 4583 7588 4639 7644
rect 4639 7588 4643 7644
rect 4579 7584 4643 7588
rect 4659 7644 4723 7648
rect 4659 7588 4663 7644
rect 4663 7588 4719 7644
rect 4719 7588 4723 7644
rect 4659 7584 4723 7588
rect 4739 7644 4803 7648
rect 4739 7588 4743 7644
rect 4743 7588 4799 7644
rect 4799 7588 4803 7644
rect 4739 7584 4803 7588
rect 4819 7644 4883 7648
rect 4819 7588 4823 7644
rect 4823 7588 4879 7644
rect 4879 7588 4883 7644
rect 4819 7584 4883 7588
rect 6557 7644 6621 7648
rect 6557 7588 6561 7644
rect 6561 7588 6617 7644
rect 6617 7588 6621 7644
rect 6557 7584 6621 7588
rect 6637 7644 6701 7648
rect 6637 7588 6641 7644
rect 6641 7588 6697 7644
rect 6697 7588 6701 7644
rect 6637 7584 6701 7588
rect 6717 7644 6781 7648
rect 6717 7588 6721 7644
rect 6721 7588 6777 7644
rect 6777 7588 6781 7644
rect 6717 7584 6781 7588
rect 6797 7644 6861 7648
rect 6797 7588 6801 7644
rect 6801 7588 6857 7644
rect 6857 7588 6861 7644
rect 6797 7584 6861 7588
rect 8535 7644 8599 7648
rect 8535 7588 8539 7644
rect 8539 7588 8595 7644
rect 8595 7588 8599 7644
rect 8535 7584 8599 7588
rect 8615 7644 8679 7648
rect 8615 7588 8619 7644
rect 8619 7588 8675 7644
rect 8675 7588 8679 7644
rect 8615 7584 8679 7588
rect 8695 7644 8759 7648
rect 8695 7588 8699 7644
rect 8699 7588 8755 7644
rect 8755 7588 8759 7644
rect 8695 7584 8759 7588
rect 8775 7644 8839 7648
rect 8775 7588 8779 7644
rect 8779 7588 8835 7644
rect 8835 7588 8839 7644
rect 8775 7584 8839 7588
rect 1941 7100 2005 7104
rect 1941 7044 1945 7100
rect 1945 7044 2001 7100
rect 2001 7044 2005 7100
rect 1941 7040 2005 7044
rect 2021 7100 2085 7104
rect 2021 7044 2025 7100
rect 2025 7044 2081 7100
rect 2081 7044 2085 7100
rect 2021 7040 2085 7044
rect 2101 7100 2165 7104
rect 2101 7044 2105 7100
rect 2105 7044 2161 7100
rect 2161 7044 2165 7100
rect 2101 7040 2165 7044
rect 2181 7100 2245 7104
rect 2181 7044 2185 7100
rect 2185 7044 2241 7100
rect 2241 7044 2245 7100
rect 2181 7040 2245 7044
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 5897 7100 5961 7104
rect 5897 7044 5901 7100
rect 5901 7044 5957 7100
rect 5957 7044 5961 7100
rect 5897 7040 5961 7044
rect 5977 7100 6041 7104
rect 5977 7044 5981 7100
rect 5981 7044 6037 7100
rect 6037 7044 6041 7100
rect 5977 7040 6041 7044
rect 6057 7100 6121 7104
rect 6057 7044 6061 7100
rect 6061 7044 6117 7100
rect 6117 7044 6121 7100
rect 6057 7040 6121 7044
rect 6137 7100 6201 7104
rect 6137 7044 6141 7100
rect 6141 7044 6197 7100
rect 6197 7044 6201 7100
rect 6137 7040 6201 7044
rect 7875 7100 7939 7104
rect 7875 7044 7879 7100
rect 7879 7044 7935 7100
rect 7935 7044 7939 7100
rect 7875 7040 7939 7044
rect 7955 7100 8019 7104
rect 7955 7044 7959 7100
rect 7959 7044 8015 7100
rect 8015 7044 8019 7100
rect 7955 7040 8019 7044
rect 8035 7100 8099 7104
rect 8035 7044 8039 7100
rect 8039 7044 8095 7100
rect 8095 7044 8099 7100
rect 8035 7040 8099 7044
rect 8115 7100 8179 7104
rect 8115 7044 8119 7100
rect 8119 7044 8175 7100
rect 8175 7044 8179 7100
rect 8115 7040 8179 7044
rect 796 6836 860 6900
rect 796 6624 860 6628
rect 796 6568 846 6624
rect 846 6568 860 6624
rect 796 6564 860 6568
rect 2601 6556 2665 6560
rect 2601 6500 2605 6556
rect 2605 6500 2661 6556
rect 2661 6500 2665 6556
rect 2601 6496 2665 6500
rect 2681 6556 2745 6560
rect 2681 6500 2685 6556
rect 2685 6500 2741 6556
rect 2741 6500 2745 6556
rect 2681 6496 2745 6500
rect 2761 6556 2825 6560
rect 2761 6500 2765 6556
rect 2765 6500 2821 6556
rect 2821 6500 2825 6556
rect 2761 6496 2825 6500
rect 2841 6556 2905 6560
rect 2841 6500 2845 6556
rect 2845 6500 2901 6556
rect 2901 6500 2905 6556
rect 2841 6496 2905 6500
rect 4579 6556 4643 6560
rect 4579 6500 4583 6556
rect 4583 6500 4639 6556
rect 4639 6500 4643 6556
rect 4579 6496 4643 6500
rect 4659 6556 4723 6560
rect 4659 6500 4663 6556
rect 4663 6500 4719 6556
rect 4719 6500 4723 6556
rect 4659 6496 4723 6500
rect 4739 6556 4803 6560
rect 4739 6500 4743 6556
rect 4743 6500 4799 6556
rect 4799 6500 4803 6556
rect 4739 6496 4803 6500
rect 4819 6556 4883 6560
rect 4819 6500 4823 6556
rect 4823 6500 4879 6556
rect 4879 6500 4883 6556
rect 4819 6496 4883 6500
rect 6557 6556 6621 6560
rect 6557 6500 6561 6556
rect 6561 6500 6617 6556
rect 6617 6500 6621 6556
rect 6557 6496 6621 6500
rect 6637 6556 6701 6560
rect 6637 6500 6641 6556
rect 6641 6500 6697 6556
rect 6697 6500 6701 6556
rect 6637 6496 6701 6500
rect 6717 6556 6781 6560
rect 6717 6500 6721 6556
rect 6721 6500 6777 6556
rect 6777 6500 6781 6556
rect 6717 6496 6781 6500
rect 6797 6556 6861 6560
rect 6797 6500 6801 6556
rect 6801 6500 6857 6556
rect 6857 6500 6861 6556
rect 6797 6496 6861 6500
rect 8535 6556 8599 6560
rect 8535 6500 8539 6556
rect 8539 6500 8595 6556
rect 8595 6500 8599 6556
rect 8535 6496 8599 6500
rect 8615 6556 8679 6560
rect 8615 6500 8619 6556
rect 8619 6500 8675 6556
rect 8675 6500 8679 6556
rect 8615 6496 8679 6500
rect 8695 6556 8759 6560
rect 8695 6500 8699 6556
rect 8699 6500 8755 6556
rect 8755 6500 8759 6556
rect 8695 6496 8759 6500
rect 8775 6556 8839 6560
rect 8775 6500 8779 6556
rect 8779 6500 8835 6556
rect 8835 6500 8839 6556
rect 8775 6496 8839 6500
rect 796 6156 860 6220
rect 1941 6012 2005 6016
rect 1941 5956 1945 6012
rect 1945 5956 2001 6012
rect 2001 5956 2005 6012
rect 1941 5952 2005 5956
rect 2021 6012 2085 6016
rect 2021 5956 2025 6012
rect 2025 5956 2081 6012
rect 2081 5956 2085 6012
rect 2021 5952 2085 5956
rect 2101 6012 2165 6016
rect 2101 5956 2105 6012
rect 2105 5956 2161 6012
rect 2161 5956 2165 6012
rect 2101 5952 2165 5956
rect 2181 6012 2245 6016
rect 2181 5956 2185 6012
rect 2185 5956 2241 6012
rect 2241 5956 2245 6012
rect 2181 5952 2245 5956
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 5897 6012 5961 6016
rect 5897 5956 5901 6012
rect 5901 5956 5957 6012
rect 5957 5956 5961 6012
rect 5897 5952 5961 5956
rect 5977 6012 6041 6016
rect 5977 5956 5981 6012
rect 5981 5956 6037 6012
rect 6037 5956 6041 6012
rect 5977 5952 6041 5956
rect 6057 6012 6121 6016
rect 6057 5956 6061 6012
rect 6061 5956 6117 6012
rect 6117 5956 6121 6012
rect 6057 5952 6121 5956
rect 6137 6012 6201 6016
rect 6137 5956 6141 6012
rect 6141 5956 6197 6012
rect 6197 5956 6201 6012
rect 6137 5952 6201 5956
rect 7875 6012 7939 6016
rect 7875 5956 7879 6012
rect 7879 5956 7935 6012
rect 7935 5956 7939 6012
rect 7875 5952 7939 5956
rect 7955 6012 8019 6016
rect 7955 5956 7959 6012
rect 7959 5956 8015 6012
rect 8015 5956 8019 6012
rect 7955 5952 8019 5956
rect 8035 6012 8099 6016
rect 8035 5956 8039 6012
rect 8039 5956 8095 6012
rect 8095 5956 8099 6012
rect 8035 5952 8099 5956
rect 8115 6012 8179 6016
rect 8115 5956 8119 6012
rect 8119 5956 8175 6012
rect 8175 5956 8179 6012
rect 8115 5952 8179 5956
rect 796 5944 860 5948
rect 796 5888 846 5944
rect 846 5888 860 5944
rect 796 5884 860 5888
rect 2601 5468 2665 5472
rect 2601 5412 2605 5468
rect 2605 5412 2661 5468
rect 2661 5412 2665 5468
rect 2601 5408 2665 5412
rect 2681 5468 2745 5472
rect 2681 5412 2685 5468
rect 2685 5412 2741 5468
rect 2741 5412 2745 5468
rect 2681 5408 2745 5412
rect 2761 5468 2825 5472
rect 2761 5412 2765 5468
rect 2765 5412 2821 5468
rect 2821 5412 2825 5468
rect 2761 5408 2825 5412
rect 2841 5468 2905 5472
rect 2841 5412 2845 5468
rect 2845 5412 2901 5468
rect 2901 5412 2905 5468
rect 2841 5408 2905 5412
rect 4579 5468 4643 5472
rect 4579 5412 4583 5468
rect 4583 5412 4639 5468
rect 4639 5412 4643 5468
rect 4579 5408 4643 5412
rect 4659 5468 4723 5472
rect 4659 5412 4663 5468
rect 4663 5412 4719 5468
rect 4719 5412 4723 5468
rect 4659 5408 4723 5412
rect 4739 5468 4803 5472
rect 4739 5412 4743 5468
rect 4743 5412 4799 5468
rect 4799 5412 4803 5468
rect 4739 5408 4803 5412
rect 4819 5468 4883 5472
rect 4819 5412 4823 5468
rect 4823 5412 4879 5468
rect 4879 5412 4883 5468
rect 4819 5408 4883 5412
rect 6557 5468 6621 5472
rect 6557 5412 6561 5468
rect 6561 5412 6617 5468
rect 6617 5412 6621 5468
rect 6557 5408 6621 5412
rect 6637 5468 6701 5472
rect 6637 5412 6641 5468
rect 6641 5412 6697 5468
rect 6697 5412 6701 5468
rect 6637 5408 6701 5412
rect 6717 5468 6781 5472
rect 6717 5412 6721 5468
rect 6721 5412 6777 5468
rect 6777 5412 6781 5468
rect 6717 5408 6781 5412
rect 6797 5468 6861 5472
rect 6797 5412 6801 5468
rect 6801 5412 6857 5468
rect 6857 5412 6861 5468
rect 6797 5408 6861 5412
rect 8535 5468 8599 5472
rect 8535 5412 8539 5468
rect 8539 5412 8595 5468
rect 8595 5412 8599 5468
rect 8535 5408 8599 5412
rect 8615 5468 8679 5472
rect 8615 5412 8619 5468
rect 8619 5412 8675 5468
rect 8675 5412 8679 5468
rect 8615 5408 8679 5412
rect 8695 5468 8759 5472
rect 8695 5412 8699 5468
rect 8699 5412 8755 5468
rect 8755 5412 8759 5468
rect 8695 5408 8759 5412
rect 8775 5468 8839 5472
rect 8775 5412 8779 5468
rect 8779 5412 8835 5468
rect 8835 5412 8839 5468
rect 8775 5408 8839 5412
rect 1941 4924 2005 4928
rect 1941 4868 1945 4924
rect 1945 4868 2001 4924
rect 2001 4868 2005 4924
rect 1941 4864 2005 4868
rect 2021 4924 2085 4928
rect 2021 4868 2025 4924
rect 2025 4868 2081 4924
rect 2081 4868 2085 4924
rect 2021 4864 2085 4868
rect 2101 4924 2165 4928
rect 2101 4868 2105 4924
rect 2105 4868 2161 4924
rect 2161 4868 2165 4924
rect 2101 4864 2165 4868
rect 2181 4924 2245 4928
rect 2181 4868 2185 4924
rect 2185 4868 2241 4924
rect 2241 4868 2245 4924
rect 2181 4864 2245 4868
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 5897 4924 5961 4928
rect 5897 4868 5901 4924
rect 5901 4868 5957 4924
rect 5957 4868 5961 4924
rect 5897 4864 5961 4868
rect 5977 4924 6041 4928
rect 5977 4868 5981 4924
rect 5981 4868 6037 4924
rect 6037 4868 6041 4924
rect 5977 4864 6041 4868
rect 6057 4924 6121 4928
rect 6057 4868 6061 4924
rect 6061 4868 6117 4924
rect 6117 4868 6121 4924
rect 6057 4864 6121 4868
rect 6137 4924 6201 4928
rect 6137 4868 6141 4924
rect 6141 4868 6197 4924
rect 6197 4868 6201 4924
rect 6137 4864 6201 4868
rect 7875 4924 7939 4928
rect 7875 4868 7879 4924
rect 7879 4868 7935 4924
rect 7935 4868 7939 4924
rect 7875 4864 7939 4868
rect 7955 4924 8019 4928
rect 7955 4868 7959 4924
rect 7959 4868 8015 4924
rect 8015 4868 8019 4924
rect 7955 4864 8019 4868
rect 8035 4924 8099 4928
rect 8035 4868 8039 4924
rect 8039 4868 8095 4924
rect 8095 4868 8099 4924
rect 8035 4864 8099 4868
rect 8115 4924 8179 4928
rect 8115 4868 8119 4924
rect 8119 4868 8175 4924
rect 8175 4868 8179 4924
rect 8115 4864 8179 4868
rect 2601 4380 2665 4384
rect 2601 4324 2605 4380
rect 2605 4324 2661 4380
rect 2661 4324 2665 4380
rect 2601 4320 2665 4324
rect 2681 4380 2745 4384
rect 2681 4324 2685 4380
rect 2685 4324 2741 4380
rect 2741 4324 2745 4380
rect 2681 4320 2745 4324
rect 2761 4380 2825 4384
rect 2761 4324 2765 4380
rect 2765 4324 2821 4380
rect 2821 4324 2825 4380
rect 2761 4320 2825 4324
rect 2841 4380 2905 4384
rect 2841 4324 2845 4380
rect 2845 4324 2901 4380
rect 2901 4324 2905 4380
rect 2841 4320 2905 4324
rect 4579 4380 4643 4384
rect 4579 4324 4583 4380
rect 4583 4324 4639 4380
rect 4639 4324 4643 4380
rect 4579 4320 4643 4324
rect 4659 4380 4723 4384
rect 4659 4324 4663 4380
rect 4663 4324 4719 4380
rect 4719 4324 4723 4380
rect 4659 4320 4723 4324
rect 4739 4380 4803 4384
rect 4739 4324 4743 4380
rect 4743 4324 4799 4380
rect 4799 4324 4803 4380
rect 4739 4320 4803 4324
rect 4819 4380 4883 4384
rect 4819 4324 4823 4380
rect 4823 4324 4879 4380
rect 4879 4324 4883 4380
rect 4819 4320 4883 4324
rect 6557 4380 6621 4384
rect 6557 4324 6561 4380
rect 6561 4324 6617 4380
rect 6617 4324 6621 4380
rect 6557 4320 6621 4324
rect 6637 4380 6701 4384
rect 6637 4324 6641 4380
rect 6641 4324 6697 4380
rect 6697 4324 6701 4380
rect 6637 4320 6701 4324
rect 6717 4380 6781 4384
rect 6717 4324 6721 4380
rect 6721 4324 6777 4380
rect 6777 4324 6781 4380
rect 6717 4320 6781 4324
rect 6797 4380 6861 4384
rect 6797 4324 6801 4380
rect 6801 4324 6857 4380
rect 6857 4324 6861 4380
rect 6797 4320 6861 4324
rect 8535 4380 8599 4384
rect 8535 4324 8539 4380
rect 8539 4324 8595 4380
rect 8595 4324 8599 4380
rect 8535 4320 8599 4324
rect 8615 4380 8679 4384
rect 8615 4324 8619 4380
rect 8619 4324 8675 4380
rect 8675 4324 8679 4380
rect 8615 4320 8679 4324
rect 8695 4380 8759 4384
rect 8695 4324 8699 4380
rect 8699 4324 8755 4380
rect 8755 4324 8759 4380
rect 8695 4320 8759 4324
rect 8775 4380 8839 4384
rect 8775 4324 8779 4380
rect 8779 4324 8835 4380
rect 8835 4324 8839 4380
rect 8775 4320 8839 4324
rect 1941 3836 2005 3840
rect 1941 3780 1945 3836
rect 1945 3780 2001 3836
rect 2001 3780 2005 3836
rect 1941 3776 2005 3780
rect 2021 3836 2085 3840
rect 2021 3780 2025 3836
rect 2025 3780 2081 3836
rect 2081 3780 2085 3836
rect 2021 3776 2085 3780
rect 2101 3836 2165 3840
rect 2101 3780 2105 3836
rect 2105 3780 2161 3836
rect 2161 3780 2165 3836
rect 2101 3776 2165 3780
rect 2181 3836 2245 3840
rect 2181 3780 2185 3836
rect 2185 3780 2241 3836
rect 2241 3780 2245 3836
rect 2181 3776 2245 3780
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 5897 3836 5961 3840
rect 5897 3780 5901 3836
rect 5901 3780 5957 3836
rect 5957 3780 5961 3836
rect 5897 3776 5961 3780
rect 5977 3836 6041 3840
rect 5977 3780 5981 3836
rect 5981 3780 6037 3836
rect 6037 3780 6041 3836
rect 5977 3776 6041 3780
rect 6057 3836 6121 3840
rect 6057 3780 6061 3836
rect 6061 3780 6117 3836
rect 6117 3780 6121 3836
rect 6057 3776 6121 3780
rect 6137 3836 6201 3840
rect 6137 3780 6141 3836
rect 6141 3780 6197 3836
rect 6197 3780 6201 3836
rect 6137 3776 6201 3780
rect 7875 3836 7939 3840
rect 7875 3780 7879 3836
rect 7879 3780 7935 3836
rect 7935 3780 7939 3836
rect 7875 3776 7939 3780
rect 7955 3836 8019 3840
rect 7955 3780 7959 3836
rect 7959 3780 8015 3836
rect 8015 3780 8019 3836
rect 7955 3776 8019 3780
rect 8035 3836 8099 3840
rect 8035 3780 8039 3836
rect 8039 3780 8095 3836
rect 8095 3780 8099 3836
rect 8035 3776 8099 3780
rect 8115 3836 8179 3840
rect 8115 3780 8119 3836
rect 8119 3780 8175 3836
rect 8175 3780 8179 3836
rect 8115 3776 8179 3780
rect 2601 3292 2665 3296
rect 2601 3236 2605 3292
rect 2605 3236 2661 3292
rect 2661 3236 2665 3292
rect 2601 3232 2665 3236
rect 2681 3292 2745 3296
rect 2681 3236 2685 3292
rect 2685 3236 2741 3292
rect 2741 3236 2745 3292
rect 2681 3232 2745 3236
rect 2761 3292 2825 3296
rect 2761 3236 2765 3292
rect 2765 3236 2821 3292
rect 2821 3236 2825 3292
rect 2761 3232 2825 3236
rect 2841 3292 2905 3296
rect 2841 3236 2845 3292
rect 2845 3236 2901 3292
rect 2901 3236 2905 3292
rect 2841 3232 2905 3236
rect 4579 3292 4643 3296
rect 4579 3236 4583 3292
rect 4583 3236 4639 3292
rect 4639 3236 4643 3292
rect 4579 3232 4643 3236
rect 4659 3292 4723 3296
rect 4659 3236 4663 3292
rect 4663 3236 4719 3292
rect 4719 3236 4723 3292
rect 4659 3232 4723 3236
rect 4739 3292 4803 3296
rect 4739 3236 4743 3292
rect 4743 3236 4799 3292
rect 4799 3236 4803 3292
rect 4739 3232 4803 3236
rect 4819 3292 4883 3296
rect 4819 3236 4823 3292
rect 4823 3236 4879 3292
rect 4879 3236 4883 3292
rect 4819 3232 4883 3236
rect 6557 3292 6621 3296
rect 6557 3236 6561 3292
rect 6561 3236 6617 3292
rect 6617 3236 6621 3292
rect 6557 3232 6621 3236
rect 6637 3292 6701 3296
rect 6637 3236 6641 3292
rect 6641 3236 6697 3292
rect 6697 3236 6701 3292
rect 6637 3232 6701 3236
rect 6717 3292 6781 3296
rect 6717 3236 6721 3292
rect 6721 3236 6777 3292
rect 6777 3236 6781 3292
rect 6717 3232 6781 3236
rect 6797 3292 6861 3296
rect 6797 3236 6801 3292
rect 6801 3236 6857 3292
rect 6857 3236 6861 3292
rect 6797 3232 6861 3236
rect 8535 3292 8599 3296
rect 8535 3236 8539 3292
rect 8539 3236 8595 3292
rect 8595 3236 8599 3292
rect 8535 3232 8599 3236
rect 8615 3292 8679 3296
rect 8615 3236 8619 3292
rect 8619 3236 8675 3292
rect 8675 3236 8679 3292
rect 8615 3232 8679 3236
rect 8695 3292 8759 3296
rect 8695 3236 8699 3292
rect 8699 3236 8755 3292
rect 8755 3236 8759 3292
rect 8695 3232 8759 3236
rect 8775 3292 8839 3296
rect 8775 3236 8779 3292
rect 8779 3236 8835 3292
rect 8835 3236 8839 3292
rect 8775 3232 8839 3236
rect 1941 2748 2005 2752
rect 1941 2692 1945 2748
rect 1945 2692 2001 2748
rect 2001 2692 2005 2748
rect 1941 2688 2005 2692
rect 2021 2748 2085 2752
rect 2021 2692 2025 2748
rect 2025 2692 2081 2748
rect 2081 2692 2085 2748
rect 2021 2688 2085 2692
rect 2101 2748 2165 2752
rect 2101 2692 2105 2748
rect 2105 2692 2161 2748
rect 2161 2692 2165 2748
rect 2101 2688 2165 2692
rect 2181 2748 2245 2752
rect 2181 2692 2185 2748
rect 2185 2692 2241 2748
rect 2241 2692 2245 2748
rect 2181 2688 2245 2692
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 5897 2748 5961 2752
rect 5897 2692 5901 2748
rect 5901 2692 5957 2748
rect 5957 2692 5961 2748
rect 5897 2688 5961 2692
rect 5977 2748 6041 2752
rect 5977 2692 5981 2748
rect 5981 2692 6037 2748
rect 6037 2692 6041 2748
rect 5977 2688 6041 2692
rect 6057 2748 6121 2752
rect 6057 2692 6061 2748
rect 6061 2692 6117 2748
rect 6117 2692 6121 2748
rect 6057 2688 6121 2692
rect 6137 2748 6201 2752
rect 6137 2692 6141 2748
rect 6141 2692 6197 2748
rect 6197 2692 6201 2748
rect 6137 2688 6201 2692
rect 7875 2748 7939 2752
rect 7875 2692 7879 2748
rect 7879 2692 7935 2748
rect 7935 2692 7939 2748
rect 7875 2688 7939 2692
rect 7955 2748 8019 2752
rect 7955 2692 7959 2748
rect 7959 2692 8015 2748
rect 8015 2692 8019 2748
rect 7955 2688 8019 2692
rect 8035 2748 8099 2752
rect 8035 2692 8039 2748
rect 8039 2692 8095 2748
rect 8095 2692 8099 2748
rect 8035 2688 8099 2692
rect 8115 2748 8179 2752
rect 8115 2692 8119 2748
rect 8119 2692 8175 2748
rect 8175 2692 8179 2748
rect 8115 2688 8179 2692
rect 2601 2204 2665 2208
rect 2601 2148 2605 2204
rect 2605 2148 2661 2204
rect 2661 2148 2665 2204
rect 2601 2144 2665 2148
rect 2681 2204 2745 2208
rect 2681 2148 2685 2204
rect 2685 2148 2741 2204
rect 2741 2148 2745 2204
rect 2681 2144 2745 2148
rect 2761 2204 2825 2208
rect 2761 2148 2765 2204
rect 2765 2148 2821 2204
rect 2821 2148 2825 2204
rect 2761 2144 2825 2148
rect 2841 2204 2905 2208
rect 2841 2148 2845 2204
rect 2845 2148 2901 2204
rect 2901 2148 2905 2204
rect 2841 2144 2905 2148
rect 4579 2204 4643 2208
rect 4579 2148 4583 2204
rect 4583 2148 4639 2204
rect 4639 2148 4643 2204
rect 4579 2144 4643 2148
rect 4659 2204 4723 2208
rect 4659 2148 4663 2204
rect 4663 2148 4719 2204
rect 4719 2148 4723 2204
rect 4659 2144 4723 2148
rect 4739 2204 4803 2208
rect 4739 2148 4743 2204
rect 4743 2148 4799 2204
rect 4799 2148 4803 2204
rect 4739 2144 4803 2148
rect 4819 2204 4883 2208
rect 4819 2148 4823 2204
rect 4823 2148 4879 2204
rect 4879 2148 4883 2204
rect 4819 2144 4883 2148
rect 6557 2204 6621 2208
rect 6557 2148 6561 2204
rect 6561 2148 6617 2204
rect 6617 2148 6621 2204
rect 6557 2144 6621 2148
rect 6637 2204 6701 2208
rect 6637 2148 6641 2204
rect 6641 2148 6697 2204
rect 6697 2148 6701 2204
rect 6637 2144 6701 2148
rect 6717 2204 6781 2208
rect 6717 2148 6721 2204
rect 6721 2148 6777 2204
rect 6777 2148 6781 2204
rect 6717 2144 6781 2148
rect 6797 2204 6861 2208
rect 6797 2148 6801 2204
rect 6801 2148 6857 2204
rect 6857 2148 6861 2204
rect 6797 2144 6861 2148
rect 8535 2204 8599 2208
rect 8535 2148 8539 2204
rect 8539 2148 8595 2204
rect 8595 2148 8599 2204
rect 8535 2144 8599 2148
rect 8615 2204 8679 2208
rect 8615 2148 8619 2204
rect 8619 2148 8675 2204
rect 8675 2148 8679 2204
rect 8615 2144 8679 2148
rect 8695 2204 8759 2208
rect 8695 2148 8699 2204
rect 8699 2148 8755 2204
rect 8755 2148 8759 2204
rect 8695 2144 8759 2148
rect 8775 2204 8839 2208
rect 8775 2148 8779 2204
rect 8779 2148 8835 2204
rect 8835 2148 8839 2204
rect 8775 2144 8839 2148
<< metal4 >>
rect 1933 9280 2253 9840
rect 1933 9216 1941 9280
rect 2005 9216 2021 9280
rect 2085 9216 2101 9280
rect 2165 9216 2181 9280
rect 2245 9216 2253 9280
rect 1933 8958 2253 9216
rect 1933 8722 1975 8958
rect 2211 8722 2253 8958
rect 1933 8192 2253 8722
rect 1933 8128 1941 8192
rect 2005 8128 2021 8192
rect 2085 8128 2101 8192
rect 2165 8128 2181 8192
rect 2245 8128 2253 8192
rect 1933 7104 2253 8128
rect 1933 7040 1941 7104
rect 2005 7054 2021 7104
rect 2085 7054 2101 7104
rect 2165 7054 2181 7104
rect 2245 7040 2253 7104
rect 795 6900 861 6901
rect 795 6836 796 6900
rect 860 6836 861 6900
rect 795 6835 861 6836
rect 798 6629 858 6835
rect 1933 6818 1975 7040
rect 2211 6818 2253 7040
rect 795 6628 861 6629
rect 795 6564 796 6628
rect 860 6564 861 6628
rect 795 6563 861 6564
rect 795 6220 861 6221
rect 795 6156 796 6220
rect 860 6156 861 6220
rect 795 6155 861 6156
rect 798 5949 858 6155
rect 1933 6016 2253 6818
rect 1933 5952 1941 6016
rect 2005 5952 2021 6016
rect 2085 5952 2101 6016
rect 2165 5952 2181 6016
rect 2245 5952 2253 6016
rect 795 5948 861 5949
rect 795 5884 796 5948
rect 860 5884 861 5948
rect 795 5883 861 5884
rect 1933 5150 2253 5952
rect 1933 4928 1975 5150
rect 2211 4928 2253 5150
rect 1933 4864 1941 4928
rect 2005 4864 2021 4914
rect 2085 4864 2101 4914
rect 2165 4864 2181 4914
rect 2245 4864 2253 4928
rect 1933 3840 2253 4864
rect 1933 3776 1941 3840
rect 2005 3776 2021 3840
rect 2085 3776 2101 3840
rect 2165 3776 2181 3840
rect 2245 3776 2253 3840
rect 1933 3246 2253 3776
rect 1933 3010 1975 3246
rect 2211 3010 2253 3246
rect 1933 2752 2253 3010
rect 1933 2688 1941 2752
rect 2005 2688 2021 2752
rect 2085 2688 2101 2752
rect 2165 2688 2181 2752
rect 2245 2688 2253 2752
rect 1933 2128 2253 2688
rect 2593 9824 2913 9840
rect 2593 9760 2601 9824
rect 2665 9760 2681 9824
rect 2745 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2913 9824
rect 2593 9618 2913 9760
rect 2593 9382 2635 9618
rect 2871 9382 2913 9618
rect 2593 8736 2913 9382
rect 2593 8672 2601 8736
rect 2665 8672 2681 8736
rect 2745 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2913 8736
rect 2593 7714 2913 8672
rect 2593 7648 2635 7714
rect 2871 7648 2913 7714
rect 2593 7584 2601 7648
rect 2905 7584 2913 7648
rect 2593 7478 2635 7584
rect 2871 7478 2913 7584
rect 2593 6560 2913 7478
rect 2593 6496 2601 6560
rect 2665 6496 2681 6560
rect 2745 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2913 6560
rect 2593 5810 2913 6496
rect 2593 5574 2635 5810
rect 2871 5574 2913 5810
rect 2593 5472 2913 5574
rect 2593 5408 2601 5472
rect 2665 5408 2681 5472
rect 2745 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2913 5472
rect 2593 4384 2913 5408
rect 2593 4320 2601 4384
rect 2665 4320 2681 4384
rect 2745 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2913 4384
rect 2593 3906 2913 4320
rect 2593 3670 2635 3906
rect 2871 3670 2913 3906
rect 2593 3296 2913 3670
rect 2593 3232 2601 3296
rect 2665 3232 2681 3296
rect 2745 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2913 3296
rect 2593 2208 2913 3232
rect 2593 2144 2601 2208
rect 2665 2144 2681 2208
rect 2745 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2913 2208
rect 2593 2128 2913 2144
rect 3911 9280 4231 9840
rect 3911 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4231 9280
rect 3911 8958 4231 9216
rect 3911 8722 3953 8958
rect 4189 8722 4231 8958
rect 3911 8192 4231 8722
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7054 3999 7104
rect 4063 7054 4079 7104
rect 4143 7054 4159 7104
rect 4223 7040 4231 7104
rect 3911 6818 3953 7040
rect 4189 6818 4231 7040
rect 3911 6016 4231 6818
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 5150 4231 5952
rect 3911 4928 3953 5150
rect 4189 4928 4231 5150
rect 3911 4864 3919 4928
rect 3983 4864 3999 4914
rect 4063 4864 4079 4914
rect 4143 4864 4159 4914
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 3246 4231 3776
rect 3911 3010 3953 3246
rect 4189 3010 4231 3246
rect 3911 2752 4231 3010
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 2128 4231 2688
rect 4571 9824 4891 9840
rect 4571 9760 4579 9824
rect 4643 9760 4659 9824
rect 4723 9760 4739 9824
rect 4803 9760 4819 9824
rect 4883 9760 4891 9824
rect 4571 9618 4891 9760
rect 4571 9382 4613 9618
rect 4849 9382 4891 9618
rect 4571 8736 4891 9382
rect 4571 8672 4579 8736
rect 4643 8672 4659 8736
rect 4723 8672 4739 8736
rect 4803 8672 4819 8736
rect 4883 8672 4891 8736
rect 4571 7714 4891 8672
rect 4571 7648 4613 7714
rect 4849 7648 4891 7714
rect 4571 7584 4579 7648
rect 4883 7584 4891 7648
rect 4571 7478 4613 7584
rect 4849 7478 4891 7584
rect 4571 6560 4891 7478
rect 4571 6496 4579 6560
rect 4643 6496 4659 6560
rect 4723 6496 4739 6560
rect 4803 6496 4819 6560
rect 4883 6496 4891 6560
rect 4571 5810 4891 6496
rect 4571 5574 4613 5810
rect 4849 5574 4891 5810
rect 4571 5472 4891 5574
rect 4571 5408 4579 5472
rect 4643 5408 4659 5472
rect 4723 5408 4739 5472
rect 4803 5408 4819 5472
rect 4883 5408 4891 5472
rect 4571 4384 4891 5408
rect 4571 4320 4579 4384
rect 4643 4320 4659 4384
rect 4723 4320 4739 4384
rect 4803 4320 4819 4384
rect 4883 4320 4891 4384
rect 4571 3906 4891 4320
rect 4571 3670 4613 3906
rect 4849 3670 4891 3906
rect 4571 3296 4891 3670
rect 4571 3232 4579 3296
rect 4643 3232 4659 3296
rect 4723 3232 4739 3296
rect 4803 3232 4819 3296
rect 4883 3232 4891 3296
rect 4571 2208 4891 3232
rect 4571 2144 4579 2208
rect 4643 2144 4659 2208
rect 4723 2144 4739 2208
rect 4803 2144 4819 2208
rect 4883 2144 4891 2208
rect 4571 2128 4891 2144
rect 5889 9280 6209 9840
rect 5889 9216 5897 9280
rect 5961 9216 5977 9280
rect 6041 9216 6057 9280
rect 6121 9216 6137 9280
rect 6201 9216 6209 9280
rect 5889 8958 6209 9216
rect 5889 8722 5931 8958
rect 6167 8722 6209 8958
rect 5889 8192 6209 8722
rect 5889 8128 5897 8192
rect 5961 8128 5977 8192
rect 6041 8128 6057 8192
rect 6121 8128 6137 8192
rect 6201 8128 6209 8192
rect 5889 7104 6209 8128
rect 5889 7040 5897 7104
rect 5961 7054 5977 7104
rect 6041 7054 6057 7104
rect 6121 7054 6137 7104
rect 6201 7040 6209 7104
rect 5889 6818 5931 7040
rect 6167 6818 6209 7040
rect 5889 6016 6209 6818
rect 5889 5952 5897 6016
rect 5961 5952 5977 6016
rect 6041 5952 6057 6016
rect 6121 5952 6137 6016
rect 6201 5952 6209 6016
rect 5889 5150 6209 5952
rect 5889 4928 5931 5150
rect 6167 4928 6209 5150
rect 5889 4864 5897 4928
rect 5961 4864 5977 4914
rect 6041 4864 6057 4914
rect 6121 4864 6137 4914
rect 6201 4864 6209 4928
rect 5889 3840 6209 4864
rect 5889 3776 5897 3840
rect 5961 3776 5977 3840
rect 6041 3776 6057 3840
rect 6121 3776 6137 3840
rect 6201 3776 6209 3840
rect 5889 3246 6209 3776
rect 5889 3010 5931 3246
rect 6167 3010 6209 3246
rect 5889 2752 6209 3010
rect 5889 2688 5897 2752
rect 5961 2688 5977 2752
rect 6041 2688 6057 2752
rect 6121 2688 6137 2752
rect 6201 2688 6209 2752
rect 5889 2128 6209 2688
rect 6549 9824 6869 9840
rect 6549 9760 6557 9824
rect 6621 9760 6637 9824
rect 6701 9760 6717 9824
rect 6781 9760 6797 9824
rect 6861 9760 6869 9824
rect 6549 9618 6869 9760
rect 6549 9382 6591 9618
rect 6827 9382 6869 9618
rect 6549 8736 6869 9382
rect 6549 8672 6557 8736
rect 6621 8672 6637 8736
rect 6701 8672 6717 8736
rect 6781 8672 6797 8736
rect 6861 8672 6869 8736
rect 6549 7714 6869 8672
rect 6549 7648 6591 7714
rect 6827 7648 6869 7714
rect 6549 7584 6557 7648
rect 6861 7584 6869 7648
rect 6549 7478 6591 7584
rect 6827 7478 6869 7584
rect 6549 6560 6869 7478
rect 6549 6496 6557 6560
rect 6621 6496 6637 6560
rect 6701 6496 6717 6560
rect 6781 6496 6797 6560
rect 6861 6496 6869 6560
rect 6549 5810 6869 6496
rect 6549 5574 6591 5810
rect 6827 5574 6869 5810
rect 6549 5472 6869 5574
rect 6549 5408 6557 5472
rect 6621 5408 6637 5472
rect 6701 5408 6717 5472
rect 6781 5408 6797 5472
rect 6861 5408 6869 5472
rect 6549 4384 6869 5408
rect 6549 4320 6557 4384
rect 6621 4320 6637 4384
rect 6701 4320 6717 4384
rect 6781 4320 6797 4384
rect 6861 4320 6869 4384
rect 6549 3906 6869 4320
rect 6549 3670 6591 3906
rect 6827 3670 6869 3906
rect 6549 3296 6869 3670
rect 6549 3232 6557 3296
rect 6621 3232 6637 3296
rect 6701 3232 6717 3296
rect 6781 3232 6797 3296
rect 6861 3232 6869 3296
rect 6549 2208 6869 3232
rect 6549 2144 6557 2208
rect 6621 2144 6637 2208
rect 6701 2144 6717 2208
rect 6781 2144 6797 2208
rect 6861 2144 6869 2208
rect 6549 2128 6869 2144
rect 7867 9280 8187 9840
rect 7867 9216 7875 9280
rect 7939 9216 7955 9280
rect 8019 9216 8035 9280
rect 8099 9216 8115 9280
rect 8179 9216 8187 9280
rect 7867 8958 8187 9216
rect 7867 8722 7909 8958
rect 8145 8722 8187 8958
rect 7867 8192 8187 8722
rect 7867 8128 7875 8192
rect 7939 8128 7955 8192
rect 8019 8128 8035 8192
rect 8099 8128 8115 8192
rect 8179 8128 8187 8192
rect 7867 7104 8187 8128
rect 7867 7040 7875 7104
rect 7939 7054 7955 7104
rect 8019 7054 8035 7104
rect 8099 7054 8115 7104
rect 8179 7040 8187 7104
rect 7867 6818 7909 7040
rect 8145 6818 8187 7040
rect 7867 6016 8187 6818
rect 7867 5952 7875 6016
rect 7939 5952 7955 6016
rect 8019 5952 8035 6016
rect 8099 5952 8115 6016
rect 8179 5952 8187 6016
rect 7867 5150 8187 5952
rect 7867 4928 7909 5150
rect 8145 4928 8187 5150
rect 7867 4864 7875 4928
rect 7939 4864 7955 4914
rect 8019 4864 8035 4914
rect 8099 4864 8115 4914
rect 8179 4864 8187 4928
rect 7867 3840 8187 4864
rect 7867 3776 7875 3840
rect 7939 3776 7955 3840
rect 8019 3776 8035 3840
rect 8099 3776 8115 3840
rect 8179 3776 8187 3840
rect 7867 3246 8187 3776
rect 7867 3010 7909 3246
rect 8145 3010 8187 3246
rect 7867 2752 8187 3010
rect 7867 2688 7875 2752
rect 7939 2688 7955 2752
rect 8019 2688 8035 2752
rect 8099 2688 8115 2752
rect 8179 2688 8187 2752
rect 7867 2128 8187 2688
rect 8527 9824 8847 9840
rect 8527 9760 8535 9824
rect 8599 9760 8615 9824
rect 8679 9760 8695 9824
rect 8759 9760 8775 9824
rect 8839 9760 8847 9824
rect 8527 9618 8847 9760
rect 8527 9382 8569 9618
rect 8805 9382 8847 9618
rect 8527 8736 8847 9382
rect 8527 8672 8535 8736
rect 8599 8672 8615 8736
rect 8679 8672 8695 8736
rect 8759 8672 8775 8736
rect 8839 8672 8847 8736
rect 8527 7714 8847 8672
rect 8527 7648 8569 7714
rect 8805 7648 8847 7714
rect 8527 7584 8535 7648
rect 8839 7584 8847 7648
rect 8527 7478 8569 7584
rect 8805 7478 8847 7584
rect 8527 6560 8847 7478
rect 8527 6496 8535 6560
rect 8599 6496 8615 6560
rect 8679 6496 8695 6560
rect 8759 6496 8775 6560
rect 8839 6496 8847 6560
rect 8527 5810 8847 6496
rect 8527 5574 8569 5810
rect 8805 5574 8847 5810
rect 8527 5472 8847 5574
rect 8527 5408 8535 5472
rect 8599 5408 8615 5472
rect 8679 5408 8695 5472
rect 8759 5408 8775 5472
rect 8839 5408 8847 5472
rect 8527 4384 8847 5408
rect 8527 4320 8535 4384
rect 8599 4320 8615 4384
rect 8679 4320 8695 4384
rect 8759 4320 8775 4384
rect 8839 4320 8847 4384
rect 8527 3906 8847 4320
rect 8527 3670 8569 3906
rect 8805 3670 8847 3906
rect 8527 3296 8847 3670
rect 8527 3232 8535 3296
rect 8599 3232 8615 3296
rect 8679 3232 8695 3296
rect 8759 3232 8775 3296
rect 8839 3232 8847 3296
rect 8527 2208 8847 3232
rect 8527 2144 8535 2208
rect 8599 2144 8615 2208
rect 8679 2144 8695 2208
rect 8759 2144 8775 2208
rect 8839 2144 8847 2208
rect 8527 2128 8847 2144
<< via4 >>
rect 1975 8722 2211 8958
rect 1975 7040 2005 7054
rect 2005 7040 2021 7054
rect 2021 7040 2085 7054
rect 2085 7040 2101 7054
rect 2101 7040 2165 7054
rect 2165 7040 2181 7054
rect 2181 7040 2211 7054
rect 1975 6818 2211 7040
rect 1975 4928 2211 5150
rect 1975 4914 2005 4928
rect 2005 4914 2021 4928
rect 2021 4914 2085 4928
rect 2085 4914 2101 4928
rect 2101 4914 2165 4928
rect 2165 4914 2181 4928
rect 2181 4914 2211 4928
rect 1975 3010 2211 3246
rect 2635 9382 2871 9618
rect 2635 7648 2871 7714
rect 2635 7584 2665 7648
rect 2665 7584 2681 7648
rect 2681 7584 2745 7648
rect 2745 7584 2761 7648
rect 2761 7584 2825 7648
rect 2825 7584 2841 7648
rect 2841 7584 2871 7648
rect 2635 7478 2871 7584
rect 2635 5574 2871 5810
rect 2635 3670 2871 3906
rect 3953 8722 4189 8958
rect 3953 7040 3983 7054
rect 3983 7040 3999 7054
rect 3999 7040 4063 7054
rect 4063 7040 4079 7054
rect 4079 7040 4143 7054
rect 4143 7040 4159 7054
rect 4159 7040 4189 7054
rect 3953 6818 4189 7040
rect 3953 4928 4189 5150
rect 3953 4914 3983 4928
rect 3983 4914 3999 4928
rect 3999 4914 4063 4928
rect 4063 4914 4079 4928
rect 4079 4914 4143 4928
rect 4143 4914 4159 4928
rect 4159 4914 4189 4928
rect 3953 3010 4189 3246
rect 4613 9382 4849 9618
rect 4613 7648 4849 7714
rect 4613 7584 4643 7648
rect 4643 7584 4659 7648
rect 4659 7584 4723 7648
rect 4723 7584 4739 7648
rect 4739 7584 4803 7648
rect 4803 7584 4819 7648
rect 4819 7584 4849 7648
rect 4613 7478 4849 7584
rect 4613 5574 4849 5810
rect 4613 3670 4849 3906
rect 5931 8722 6167 8958
rect 5931 7040 5961 7054
rect 5961 7040 5977 7054
rect 5977 7040 6041 7054
rect 6041 7040 6057 7054
rect 6057 7040 6121 7054
rect 6121 7040 6137 7054
rect 6137 7040 6167 7054
rect 5931 6818 6167 7040
rect 5931 4928 6167 5150
rect 5931 4914 5961 4928
rect 5961 4914 5977 4928
rect 5977 4914 6041 4928
rect 6041 4914 6057 4928
rect 6057 4914 6121 4928
rect 6121 4914 6137 4928
rect 6137 4914 6167 4928
rect 5931 3010 6167 3246
rect 6591 9382 6827 9618
rect 6591 7648 6827 7714
rect 6591 7584 6621 7648
rect 6621 7584 6637 7648
rect 6637 7584 6701 7648
rect 6701 7584 6717 7648
rect 6717 7584 6781 7648
rect 6781 7584 6797 7648
rect 6797 7584 6827 7648
rect 6591 7478 6827 7584
rect 6591 5574 6827 5810
rect 6591 3670 6827 3906
rect 7909 8722 8145 8958
rect 7909 7040 7939 7054
rect 7939 7040 7955 7054
rect 7955 7040 8019 7054
rect 8019 7040 8035 7054
rect 8035 7040 8099 7054
rect 8099 7040 8115 7054
rect 8115 7040 8145 7054
rect 7909 6818 8145 7040
rect 7909 4928 8145 5150
rect 7909 4914 7939 4928
rect 7939 4914 7955 4928
rect 7955 4914 8019 4928
rect 8019 4914 8035 4928
rect 8035 4914 8099 4928
rect 8099 4914 8115 4928
rect 8115 4914 8145 4928
rect 7909 3010 8145 3246
rect 8569 9382 8805 9618
rect 8569 7648 8805 7714
rect 8569 7584 8599 7648
rect 8599 7584 8615 7648
rect 8615 7584 8679 7648
rect 8679 7584 8695 7648
rect 8695 7584 8759 7648
rect 8759 7584 8775 7648
rect 8775 7584 8805 7648
rect 8569 7478 8805 7584
rect 8569 5574 8805 5810
rect 8569 3670 8805 3906
<< metal5 >>
rect 1056 9618 9064 9660
rect 1056 9382 2635 9618
rect 2871 9382 4613 9618
rect 4849 9382 6591 9618
rect 6827 9382 8569 9618
rect 8805 9382 9064 9618
rect 1056 9340 9064 9382
rect 1056 8958 9064 9000
rect 1056 8722 1975 8958
rect 2211 8722 3953 8958
rect 4189 8722 5931 8958
rect 6167 8722 7909 8958
rect 8145 8722 9064 8958
rect 1056 8680 9064 8722
rect 1056 7714 9064 7756
rect 1056 7478 2635 7714
rect 2871 7478 4613 7714
rect 4849 7478 6591 7714
rect 6827 7478 8569 7714
rect 8805 7478 9064 7714
rect 1056 7436 9064 7478
rect 1056 7054 9064 7096
rect 1056 6818 1975 7054
rect 2211 6818 3953 7054
rect 4189 6818 5931 7054
rect 6167 6818 7909 7054
rect 8145 6818 9064 7054
rect 1056 6776 9064 6818
rect 1056 5810 9064 5852
rect 1056 5574 2635 5810
rect 2871 5574 4613 5810
rect 4849 5574 6591 5810
rect 6827 5574 8569 5810
rect 8805 5574 9064 5810
rect 1056 5532 9064 5574
rect 1056 5150 9064 5192
rect 1056 4914 1975 5150
rect 2211 4914 3953 5150
rect 4189 4914 5931 5150
rect 6167 4914 7909 5150
rect 8145 4914 9064 5150
rect 1056 4872 9064 4914
rect 1056 3906 9064 3948
rect 1056 3670 2635 3906
rect 2871 3670 4613 3906
rect 4849 3670 6591 3906
rect 6827 3670 8569 3906
rect 8805 3670 9064 3906
rect 1056 3628 9064 3670
rect 1056 3246 9064 3288
rect 1056 3010 1975 3246
rect 2211 3010 3953 3246
rect 4189 3010 5931 3246
rect 6167 3010 7909 3246
rect 8145 3010 9064 3246
rect 1056 2968 9064 3010
use sky130_fd_sc_hd__nor2_4  _105_
timestamp 0
transform -1 0 6072 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _106_
timestamp 0
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _107_
timestamp 0
transform 1 0 5796 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _108_
timestamp 0
transform 1 0 6440 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _109_
timestamp 0
transform -1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _110_
timestamp 0
transform -1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _111_
timestamp 0
transform -1 0 8740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _113_
timestamp 0
transform -1 0 6716 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _114_
timestamp 0
transform 1 0 5796 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_4  _115_
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_4  _116_
timestamp 0
transform -1 0 8740 0 -1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 0
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 0
transform -1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _119_
timestamp 0
transform 1 0 5428 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _120_
timestamp 0
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _121_
timestamp 0
transform -1 0 6164 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 0
transform -1 0 5704 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _123_
timestamp 0
transform 1 0 4968 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 0
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _125_
timestamp 0
transform 1 0 5520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _126_
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _127_
timestamp 0
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _128_
timestamp 0
transform -1 0 8372 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _129_
timestamp 0
transform 1 0 7728 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _130_
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _131_
timestamp 0
transform 1 0 8280 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _132_
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _133_
timestamp 0
transform -1 0 7912 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _134_
timestamp 0
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _135_
timestamp 0
transform -1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _136_
timestamp 0
transform -1 0 8464 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 0
transform -1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _139_
timestamp 0
transform -1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _140_
timestamp 0
transform 1 0 7268 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _141_
timestamp 0
transform 1 0 6716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 0
transform 1 0 8004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _143_
timestamp 0
transform 1 0 8004 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 0
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _145_
timestamp 0
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _146_
timestamp 0
transform 1 0 6624 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_2  _147_
timestamp 0
transform -1 0 6072 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _148_
timestamp 0
transform -1 0 5704 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _149_
timestamp 0
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _150_
timestamp 0
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _151_
timestamp 0
transform 1 0 6072 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _152_
timestamp 0
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 0
transform 1 0 4508 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _154_
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _155_
timestamp 0
transform -1 0 6992 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _156_
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _157_
timestamp 0
transform -1 0 4876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _158_
timestamp 0
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _159_
timestamp 0
transform 1 0 2576 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _160_
timestamp 0
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _161_
timestamp 0
transform -1 0 2392 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _162_
timestamp 0
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _163_
timestamp 0
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _164_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _165_
timestamp 0
transform 1 0 2024 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _166_
timestamp 0
transform -1 0 2024 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _167_
timestamp 0
transform -1 0 2300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 0
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _169_
timestamp 0
transform -1 0 3680 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _170_
timestamp 0
transform -1 0 4416 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 0
transform 1 0 2668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _172_
timestamp 0
transform -1 0 4600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _176_
timestamp 0
transform -1 0 2576 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _177_
timestamp 0
transform -1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _178_
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _179_
timestamp 0
transform 1 0 3036 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _180_
timestamp 0
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _181_
timestamp 0
transform -1 0 2024 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _182_
timestamp 0
transform -1 0 2392 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 0
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _184_
timestamp 0
transform 1 0 3128 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _185_
timestamp 0
transform -1 0 4784 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _186_
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _187_
timestamp 0
transform 1 0 2024 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _188_
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _189_
timestamp 0
transform 1 0 1564 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _190_
timestamp 0
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 0
transform -1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _192_
timestamp 0
transform 1 0 2392 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _193_
timestamp 0
transform 1 0 2024 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _194_
timestamp 0
transform -1 0 2024 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _195_
timestamp 0
transform -1 0 2300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 0
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _197_
timestamp 0
transform 1 0 3128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _198_
timestamp 0
transform -1 0 3128 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _199_
timestamp 0
transform 1 0 2668 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _200_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _201_
timestamp 0
transform 1 0 3772 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _202_
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _203_
timestamp 0
transform 1 0 4232 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _204_
timestamp 0
transform -1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _205_
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _206_
timestamp 0
transform 1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _207_
timestamp 0
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _208_
timestamp 0
transform -1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _209_
timestamp 0
transform 1 0 4784 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _210_
timestamp 0
transform 1 0 5520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 0
transform 1 0 3956 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _212_
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _213_
timestamp 0
transform 1 0 5060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _214_
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _215_
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _216_
timestamp 0
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 0
transform -1 0 6624 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _218_
timestamp 0
transform 1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 0
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 0
transform -1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 0
transform -1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 0
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 0
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 0
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_13
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_28
timestamp 0
transform 1 0 3680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_82
timestamp 0
transform 1 0 8648 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_13
timestamp 0
transform 1 0 2300 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_60
timestamp 0
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_13
timestamp 0
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_22
timestamp 0
transform 1 0 3128 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_28
timestamp 0
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_38
timestamp 0
transform 1 0 4600 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_82
timestamp 0
transform 1 0 8648 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_13
timestamp 0
transform 1 0 2300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_21
timestamp 0
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_29
timestamp 0
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_42
timestamp 0
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_60
timestamp 0
transform 1 0 6624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_17
timestamp 0
transform 1 0 2668 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_55
timestamp 0
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_72
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_35
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_10
timestamp 0
transform 1 0 2024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_16
timestamp 0
transform 1 0 2576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_22
timestamp 0
transform 1 0 3128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_40
timestamp 0
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_69
timestamp 0
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_13
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_25
timestamp 0
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_42
timestamp 0
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_54
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_62
timestamp 0
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_7
timestamp 0
transform 1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_16
timestamp 0
transform 1 0 2576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_28
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_36
timestamp 0
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_41
timestamp 0
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_67
timestamp 0
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_74
timestamp 0
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_82
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_14
timestamp 0
transform 1 0 2392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_59
timestamp 0
transform 1 0 6532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_82
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_6
timestamp 0
transform 1 0 1656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_13
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_29
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_67
timestamp 0
transform 1 0 7268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_78
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform -1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform -1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform -1 0 7268 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform -1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform -1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform 1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 0
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform -1 0 3680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 0
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input19
timestamp 0
transform -1 0 8740 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input20
timestamp 0
transform -1 0 8740 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output21
timestamp 0
transform -1 0 5612 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 0
transform -1 0 6256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 0
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 0
transform -1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 0
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 0
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 0
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output29
timestamp 0
transform 1 0 3956 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 9016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 9016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 9016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 9016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer1
timestamp 0
transform -1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 0
transform -1 0 3680 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 0
transform 1 0 5520 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer4
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer5
timestamp 0
transform 1 0 7268 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer6
timestamp 0
transform -1 0 8280 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 0
transform 1 0 6624 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer8
timestamp 0
transform 1 0 8004 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 0
transform -1 0 7728 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer10
timestamp 0
transform -1 0 7360 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer11
timestamp 0
transform -1 0 8004 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer12
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer13
timestamp 0
transform -1 0 4784 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_32
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_33
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_34
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_35
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_36
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_37
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_38
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_39
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_40
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_41
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_42
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_43
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
rlabel metal1 s 5060 9792 5060 9792 4 VGND
rlabel metal1 s 5060 9248 5060 9248 4 VPWR
rlabel metal1 s 2622 5746 2622 5746 4 _000_
rlabel metal1 s 2070 5712 2070 5712 4 _001_
rlabel metal1 s 2162 5712 2162 5712 4 _002_
rlabel metal1 s 2346 6324 2346 6324 4 _003_
rlabel metal1 s 3496 6222 3496 6222 4 _004_
rlabel metal2 s 1817 5610 1817 5610 4 _005_
rlabel metal2 s 1702 5916 1702 5916 4 _006_
rlabel metal2 s 3450 5372 3450 5372 4 _007_
rlabel metal1 s 2254 2278 2254 2278 4 _008_
rlabel metal1 s 4232 6290 4232 6290 4 _009_
rlabel metal1 s 2714 4148 2714 4148 4 _010_
rlabel metal2 s 1702 3162 1702 3162 4 _011_
rlabel metal1 s 1794 2618 1794 2618 4 _012_
rlabel metal1 s 1932 3162 1932 3162 4 _013_
rlabel metal1 s 1840 3706 1840 3706 4 _014_
rlabel metal1 s 2208 4522 2208 4522 4 _015_
rlabel metal1 s 2898 3706 2898 3706 4 _016_
rlabel metal1 s 1919 4182 1919 4182 4 _017_
rlabel metal2 s 1610 4284 1610 4284 4 _018_
rlabel metal1 s 2806 3060 2806 3060 4 _019_
rlabel metal1 s 3036 3026 3036 3026 4 _020_
rlabel metal2 s 4002 3264 4002 3264 4 _021_
rlabel metal1 s 3312 3978 3312 3978 4 _022_
rlabel metal1 s 3956 3434 3956 3434 4 _023_
rlabel metal1 s 4324 3162 4324 3162 4 _024_
rlabel metal1 s 3910 2618 3910 2618 4 _025_
rlabel metal1 s 5106 3094 5106 3094 4 _026_
rlabel metal1 s 5014 4012 5014 4012 4 _027_
rlabel metal2 s 4194 3434 4194 3434 4 _028_
rlabel metal1 s 4922 3570 4922 3570 4 _029_
rlabel metal2 s 4278 5474 4278 5474 4 _030_
rlabel metal1 s 5336 4114 5336 4114 4 _031_
rlabel metal2 s 5566 3196 5566 3196 4 _032_
rlabel metal1 s 5152 3570 5152 3570 4 _033_
rlabel metal2 s 5106 3264 5106 3264 4 _034_
rlabel metal1 s 7176 2822 7176 2822 4 _035_
rlabel metal1 s 6256 3434 6256 3434 4 _036_
rlabel metal1 s 4232 2550 4232 2550 4 _037_
rlabel metal1 s 6762 3638 6762 3638 4 _038_
rlabel metal2 s 1932 5610 1932 5610 4 _039_
rlabel metal1 s 6532 3026 6532 3026 4 _040_
rlabel metal2 s 6854 2346 6854 2346 4 _041_
rlabel metal1 s 7360 2414 7360 2414 4 _042_
rlabel metal2 s 2530 3196 2530 3196 4 _043_
rlabel metal1 s 7636 2618 7636 2618 4 _044_
rlabel metal1 s 8464 2618 8464 2618 4 _045_
rlabel metal1 s 2208 6290 2208 6290 4 _046_
rlabel metal1 s 6026 4624 6026 4624 4 _047_
rlabel metal2 s 6302 5440 6302 5440 4 _048_
rlabel metal2 s 7314 4590 7314 4590 4 _049_
rlabel metal2 s 7406 4590 7406 4590 4 _050_
rlabel metal3 s 5750 5219 5750 5219 4 _051_
rlabel metal1 s 6026 4250 6026 4250 4 _052_
rlabel metal1 s 1610 6358 1610 6358 4 _053_
rlabel metal1 s 7084 4250 7084 4250 4 _054_
rlabel metal2 s 6003 5270 6003 5270 4 _055_
rlabel metal1 s 7268 5746 7268 5746 4 _056_
rlabel metal2 s 6532 6290 6532 6290 4 _057_
rlabel metal1 s 6210 6290 6210 6290 4 _058_
rlabel metal2 s 6946 5474 6946 5474 4 _059_
rlabel metal1 s 6164 5202 6164 5202 4 _060_
rlabel metal1 s 8234 3162 8234 3162 4 _061_
rlabel metal1 s 8188 6766 8188 6766 4 _062_
rlabel metal2 s 7590 5474 7590 5474 4 _063_
rlabel metal1 s 8832 6698 8832 6698 4 _064_
rlabel metal1 s 7498 7854 7498 7854 4 _065_
rlabel metal2 s 7498 8092 7498 8092 4 _066_
rlabel metal1 s 8188 7718 8188 7718 4 _067_
rlabel metal1 s 8694 5644 8694 5644 4 _068_
rlabel metal1 s 8464 5678 8464 5678 4 _069_
rlabel metal1 s 7958 5882 7958 5882 4 _070_
rlabel metal1 s 7406 7412 7406 7412 4 _071_
rlabel metal2 s 7774 7718 7774 7718 4 _072_
rlabel metal2 s 7314 7344 7314 7344 4 _073_
rlabel metal1 s 8418 8466 8418 8466 4 _074_
rlabel metal1 s 7866 8602 7866 8602 4 _075_
rlabel metal2 s 8431 8942 8431 8942 4 _076_
rlabel metal1 s 7314 8908 7314 8908 4 _077_
rlabel metal1 s 5106 8942 5106 8942 4 _078_
rlabel metal1 s 5428 9486 5428 9486 4 _079_
rlabel metal2 s 4922 8092 4922 8092 4 _080_
rlabel metal1 s 4830 7888 4830 7888 4 _081_
rlabel metal2 s 5198 8840 5198 8840 4 _082_
rlabel metal2 s 6210 8636 6210 8636 4 _083_
rlabel metal1 s 5267 7786 5267 7786 4 _084_
rlabel metal1 s 5106 7514 5106 7514 4 _085_
rlabel metal1 s 5980 9554 5980 9554 4 _086_
rlabel metal1 s 3588 9146 3588 9146 4 _087_
rlabel metal2 s 6026 8636 6026 8636 4 _088_
rlabel metal2 s 2906 8602 2906 8602 4 _089_
rlabel metal1 s 3266 9078 3266 9078 4 _090_
rlabel metal1 s 2346 8908 2346 8908 4 _091_
rlabel metal1 s 1932 7446 1932 7446 4 _092_
rlabel metal1 s 2070 7344 2070 7344 4 _093_
rlabel metal2 s 2346 8092 2346 8092 4 _094_
rlabel metal1 s 4554 7820 4554 7820 4 _095_
rlabel metal2 s 1725 7446 1725 7446 4 _096_
rlabel metal2 s 1610 7548 1610 7548 4 _097_
rlabel metal1 s 4186 8500 4186 8500 4 _098_
rlabel metal1 s 4094 8432 4094 8432 4 _099_
rlabel metal1 s 4462 6970 4462 6970 4 _100_
rlabel metal1 s 3542 7922 3542 7922 4 _101_
rlabel metal2 s 4278 7242 4278 7242 4 _102_
rlabel metal1 s 3772 5882 3772 5882 4 _103_
rlabel metal2 s 3818 6154 3818 6154 4 _104_
rlabel metal1 s 2852 2414 2852 2414 4 a[0]
rlabel metal2 s 7038 3825 7038 3825 4 a[1]
rlabel metal1 s 8832 9554 8832 9554 4 a[2]
rlabel metal1 s 7222 9588 7222 9588 4 a[3]
rlabel metal3 s 866 9588 866 9588 4 a[4]
rlabel metal3 s 1004 7548 1004 7548 4 a[5]
rlabel metal2 s 2622 1027 2622 1027 4 a[6]
rlabel metal1 s 3312 3502 3312 3502 4 a[7]
rlabel metal1 s 7314 2618 7314 2618 4 alu0.result
rlabel metal1 s 5336 5202 5336 5202 4 alu1.result
rlabel metal1 s 5290 6324 5290 6324 4 alu2.result
rlabel metal2 s 4646 8262 4646 8262 4 alu3.result
rlabel metal1 s 2346 7514 2346 7514 4 alu4.result
rlabel metal2 s 2346 5916 2346 5916 4 alu5.result
rlabel metal1 s 2300 4250 2300 4250 4 alu6.result
rlabel metal1 s 4646 4250 4646 4250 4 alu7.result
rlabel metal2 s 5658 3910 5658 3910 4 b[0]
rlabel metal2 s 6210 4403 6210 4403 4 b[1]
rlabel metal2 s 7038 8381 7038 8381 4 b[2]
rlabel metal1 s 4370 9554 4370 9554 4 b[3]
rlabel metal3 s 1050 8908 1050 8908 4 b[4]
rlabel metal3 s 820 5508 820 5508 4 b[5]
rlabel metal3 s 1050 3468 1050 3468 4 b[6]
rlabel metal2 s 3910 959 3910 959 4 b[7]
rlabel metal2 s 1702 2465 1702 2465 4 cin
rlabel metal2 s 5198 1554 5198 1554 4 cout
rlabel metal1 s 3082 2346 3082 2346 4 net1
rlabel metal2 s 6394 5440 6394 5440 4 net10
rlabel metal1 s 7820 8466 7820 8466 4 net11
rlabel metal1 s 5106 9520 5106 9520 4 net12
rlabel metal1 s 3450 9554 3450 9554 4 net13
rlabel metal2 s 2438 5508 2438 5508 4 net14
rlabel metal1 s 2346 3502 2346 3502 4 net15
rlabel metal1 s 3266 3366 3266 3366 4 net16
rlabel metal2 s 1886 2108 1886 2108 4 net17
rlabel metal1 s 4462 6256 4462 6256 4 net18
rlabel metal1 s 6440 6766 6440 6766 4 net19
rlabel metal1 s 7130 5202 7130 5202 4 net2
rlabel metal1 s 7774 7854 7774 7854 4 net20
rlabel metal1 s 5612 2414 5612 2414 4 net21
rlabel metal1 s 6210 3060 6210 3060 4 net22
rlabel metal2 s 8418 4556 8418 4556 4 net23
rlabel metal1 s 5566 6154 5566 6154 4 net24
rlabel metal1 s 4922 8602 4922 8602 4 net25
rlabel metal2 s 1702 8908 1702 8908 4 net26
rlabel metal1 s 1748 6766 1748 6766 4 net27
rlabel metal1 s 1702 5168 1702 5168 4 net28
rlabel metal1 s 3910 2414 3910 2414 4 net29
rlabel metal1 s 7636 9554 7636 9554 4 net3
rlabel metal2 s 3634 9180 3634 9180 4 net30
rlabel metal1 s 2806 8466 2806 8466 4 net31
rlabel metal2 s 5658 8942 5658 8942 4 net32
rlabel metal1 s 5934 8500 5934 8500 4 net33
rlabel metal1 s 7958 5746 7958 5746 4 net34
rlabel metal1 s 7360 6902 7360 6902 4 net35
rlabel metal1 s 7866 4658 7866 4658 4 net36
rlabel metal1 s 8418 4794 8418 4794 4 net37
rlabel metal1 s 7268 4658 7268 4658 4 net38
rlabel metal2 s 6762 4998 6762 4998 4 net39
rlabel metal2 s 5566 8738 5566 8738 4 net4
rlabel metal1 s 5750 4692 5750 4692 4 net40
rlabel metal2 s 5290 4216 5290 4216 4 net41
rlabel metal2 s 4278 4454 4278 4454 4 net42
rlabel metal2 s 2622 9112 2622 9112 4 net5
rlabel metal1 s 3128 6698 3128 6698 4 net6
rlabel metal2 s 1794 2346 1794 2346 4 net7
rlabel metal1 s 3174 3604 3174 3604 4 net8
rlabel metal1 s 6118 2550 6118 2550 4 net9
rlabel metal3 s 0 6128 800 6248 4 op[0]
port 21 nsew
rlabel metal2 s 8602 6239 8602 6239 4 op[1]
rlabel metal2 s 8602 7123 8602 7123 4 op[2]
rlabel metal1 s 6256 2822 6256 2822 4 result[0]
rlabel metal1 s 8786 3978 8786 3978 4 result[1]
rlabel metal1 s 8786 7718 8786 7718 4 result[2]
rlabel metal1 s 4416 9622 4416 9622 4 result[3]
rlabel metal3 s 1096 8228 1096 8228 4 result[4]
rlabel metal3 s 0 6808 800 6928 4 result[5]
port 29 nsew
rlabel metal3 s 1096 4828 1096 4828 4 result[6]
rlabel metal2 s 4554 959 4554 959 4 result[7]
flabel metal5 s 1056 9340 9064 9660 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 7436 9064 7756 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5532 9064 5852 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3628 9064 3948 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 8527 2128 8847 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 6549 2128 6869 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4571 2128 4891 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2593 2128 2913 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8680 9064 9000 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 6776 9064 7096 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4872 9064 5192 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2968 9064 3288 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 7867 2128 8187 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5889 2128 6209 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3911 2128 4231 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1933 2128 2253 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 9401 2048 10201 2168 0 FreeSans 600 0 0 0 a[0]
port 3 nsew
flabel metal3 s 9401 4088 10201 4208 0 FreeSans 600 0 0 0 a[1]
port 4 nsew
flabel metal3 s 9401 8168 10201 8288 0 FreeSans 600 0 0 0 a[2]
port 5 nsew
flabel metal2 s 5814 11545 5870 12345 0 FreeSans 280 90 0 0 a[3]
port 6 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 a[4]
port 7 nsew
flabel metal3 s 0 7488 800 7608 0 FreeSans 600 0 0 0 a[5]
port 8 nsew
flabel metal2 s 2594 0 2650 800 0 FreeSans 280 90 0 0 a[6]
port 9 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 a[7]
port 10 nsew
flabel metal3 s 9401 3408 10201 3528 0 FreeSans 600 0 0 0 b[0]
port 11 nsew
flabel metal3 s 9401 4768 10201 4888 0 FreeSans 600 0 0 0 b[1]
port 12 nsew
flabel metal3 s 9401 8848 10201 8968 0 FreeSans 600 0 0 0 b[2]
port 13 nsew
flabel metal2 s 5170 11545 5226 12345 0 FreeSans 280 90 0 0 b[3]
port 14 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 b[4]
port 15 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 b[5]
port 16 nsew
flabel metal3 s 0 3408 800 3528 0 FreeSans 600 0 0 0 b[6]
port 17 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 b[7]
port 18 nsew
flabel metal3 s 9401 2728 10201 2848 0 FreeSans 600 0 0 0 cin
port 19 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 cout
port 20 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 op[0]
flabel metal3 s 9401 6128 10201 6248 0 FreeSans 600 0 0 0 op[1]
port 22 nsew
flabel metal3 s 9401 6808 10201 6928 0 FreeSans 600 0 0 0 op[2]
port 23 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 result[0]
port 24 nsew
flabel metal3 s 9401 5448 10201 5568 0 FreeSans 600 0 0 0 result[1]
port 25 nsew
flabel metal3 s 9401 7488 10201 7608 0 FreeSans 600 0 0 0 result[2]
port 26 nsew
flabel metal2 s 4526 11545 4582 12345 0 FreeSans 280 90 0 0 result[3]
port 27 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 result[4]
port 28 nsew
flabel metal3 s 400 6868 400 6868 0 FreeSans 600 0 0 0 result[5]
flabel metal3 s 0 4768 800 4888 0 FreeSans 600 0 0 0 result[6]
port 30 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 result[7]
port 31 nsew
<< properties >>
string FIXED_BBOX 0 0 10201 12345
<< end >>
