magic
tech sky130A
magscale 1 2
timestamp 1746639542
<< nwell >>
rect 1066 2159 9054 9809
<< obsli1 >>
rect 1104 2159 9016 9809
<< obsm1 >>
rect 842 1912 9186 9840
<< metal2 >>
rect 4526 11545 4582 12345
rect 5170 11545 5226 12345
rect 5814 11545 5870 12345
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
<< obsm2 >>
rect 846 11489 4470 11545
rect 4638 11489 5114 11545
rect 5282 11489 5758 11545
rect 5926 11489 9182 11545
rect 846 856 9182 11489
rect 846 800 2538 856
rect 2706 800 3182 856
rect 3350 800 3826 856
rect 3994 800 4470 856
rect 4638 800 5114 856
rect 5282 800 6402 856
rect 6570 800 9182 856
<< metal3 >>
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 9401 8848 10201 8968
rect 0 8168 800 8288
rect 9401 8168 10201 8288
rect 0 7488 800 7608
rect 9401 7488 10201 7608
rect 0 6808 800 6928
rect 9401 6808 10201 6928
rect 0 6128 800 6248
rect 9401 6128 10201 6248
rect 0 5448 800 5568
rect 9401 5448 10201 5568
rect 0 4768 800 4888
rect 9401 4768 10201 4888
rect 9401 4088 10201 4208
rect 0 3408 800 3528
rect 9401 3408 10201 3528
rect 9401 2728 10201 2848
rect 9401 2048 10201 2168
<< obsm3 >>
rect 750 9728 9401 9825
rect 880 9448 9401 9728
rect 750 9048 9401 9448
rect 880 8768 9321 9048
rect 750 8368 9401 8768
rect 880 8088 9321 8368
rect 750 7688 9401 8088
rect 880 7408 9321 7688
rect 750 7008 9401 7408
rect 880 6728 9321 7008
rect 750 6328 9401 6728
rect 880 6048 9321 6328
rect 750 5648 9401 6048
rect 880 5368 9321 5648
rect 750 4968 9401 5368
rect 880 4688 9321 4968
rect 750 4288 9401 4688
rect 750 4008 9321 4288
rect 750 3608 9401 4008
rect 880 3328 9321 3608
rect 750 2928 9401 3328
rect 750 2648 9321 2928
rect 750 2248 9401 2648
rect 750 1968 9321 2248
rect 750 1939 9401 1968
<< metal4 >>
rect 1933 2128 2253 9840
rect 2593 2128 2913 9840
rect 3911 2128 4231 9840
rect 4571 2128 4891 9840
rect 5889 2128 6209 9840
rect 6549 2128 6869 9840
rect 7867 2128 8187 9840
rect 8527 2128 8847 9840
<< obsm4 >>
rect 795 5883 861 6901
<< metal5 >>
rect 1056 9340 9064 9660
rect 1056 8680 9064 9000
rect 1056 7436 9064 7756
rect 1056 6776 9064 7096
rect 1056 5532 9064 5852
rect 1056 4872 9064 5192
rect 1056 3628 9064 3948
rect 1056 2968 9064 3288
<< labels >>
rlabel metal4 s 2593 2128 2913 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4571 2128 4891 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6549 2128 6869 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8527 2128 8847 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3628 9064 3948 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5532 9064 5852 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7436 9064 7756 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9340 9064 9660 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1933 2128 2253 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3911 2128 4231 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5889 2128 6209 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7867 2128 8187 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2968 9064 3288 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4872 9064 5192 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6776 9064 7096 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8680 9064 9000 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 9401 2048 10201 2168 6 a[0]
port 3 nsew signal input
rlabel metal3 s 9401 4088 10201 4208 6 a[1]
port 4 nsew signal input
rlabel metal3 s 9401 8168 10201 8288 6 a[2]
port 5 nsew signal input
rlabel metal2 s 5814 11545 5870 12345 6 a[3]
port 6 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 a[4]
port 7 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 a[5]
port 8 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 a[6]
port 9 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 a[7]
port 10 nsew signal input
rlabel metal3 s 9401 3408 10201 3528 6 b[0]
port 11 nsew signal input
rlabel metal3 s 9401 4768 10201 4888 6 b[1]
port 12 nsew signal input
rlabel metal3 s 9401 8848 10201 8968 6 b[2]
port 13 nsew signal input
rlabel metal2 s 5170 11545 5226 12345 6 b[3]
port 14 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 b[4]
port 15 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 b[5]
port 16 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 b[6]
port 17 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 b[7]
port 18 nsew signal input
rlabel metal3 s 9401 2728 10201 2848 6 cin
port 19 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 cout
port 20 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 op[0]
port 21 nsew signal input
rlabel metal3 s 9401 6128 10201 6248 6 op[1]
port 22 nsew signal input
rlabel metal3 s 9401 6808 10201 6928 6 op[2]
port 23 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 result[0]
port 24 nsew signal output
rlabel metal3 s 9401 5448 10201 5568 6 result[1]
port 25 nsew signal output
rlabel metal3 s 9401 7488 10201 7608 6 result[2]
port 26 nsew signal output
rlabel metal2 s 4526 11545 4582 12345 6 result[3]
port 27 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 result[4]
port 28 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 result[5]
port 29 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 result[6]
port 30 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 result[7]
port 31 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 10201 12345
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 724928
string GDS_FILE /openlane/designs/alu_8bit/runs/RUN_2025.05.07_17.36.09/results/signoff/alu_8bit.magic.gds
string GDS_START 312388
<< end >>

