magic
tech sky130A
magscale 1 2
timestamp 1746638556
<< nwell >>
rect 1066 2159 10894 11462
<< obsli1 >>
rect 1104 2159 10856 11441
<< obsm1 >>
rect 842 2128 10856 11892
<< metal2 >>
rect 3882 13342 3938 14142
rect 4526 13342 4582 14142
rect 5814 13342 5870 14142
rect 7102 13342 7158 14142
rect 7746 13342 7802 14142
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
<< obsm2 >>
rect 846 13286 3826 13410
rect 3994 13286 4470 13410
rect 4638 13286 5758 13410
rect 5926 13286 7046 13410
rect 7214 13286 7690 13410
rect 7858 13286 10746 13410
rect 846 856 10746 13286
rect 846 800 3826 856
rect 3994 800 4470 856
rect 4638 800 5114 856
rect 5282 800 6402 856
rect 6570 800 7046 856
rect 7214 800 7690 856
rect 7858 800 8334 856
rect 8502 800 8978 856
rect 9146 800 9622 856
rect 9790 800 10746 856
<< metal3 >>
rect 0 10208 800 10328
rect 0 8848 800 8968
rect 11198 8848 11998 8968
rect 0 8168 800 8288
rect 11198 8168 11998 8288
rect 0 7488 800 7608
rect 11198 7488 11998 7608
rect 11198 6808 11998 6928
rect 0 6128 800 6248
rect 11198 6128 11998 6248
rect 0 5448 800 5568
rect 11198 5448 11998 5568
rect 0 4768 800 4888
rect 11198 4768 11998 4888
rect 0 3408 800 3528
<< obsm3 >>
rect 798 10408 11198 11457
rect 880 10128 11198 10408
rect 798 9048 11198 10128
rect 880 8768 11118 9048
rect 798 8368 11198 8768
rect 880 8088 11118 8368
rect 798 7688 11198 8088
rect 880 7408 11118 7688
rect 798 7008 11198 7408
rect 798 6728 11118 7008
rect 798 6328 11198 6728
rect 880 6048 11118 6328
rect 798 5648 11198 6048
rect 880 5368 11118 5648
rect 798 4968 11198 5368
rect 880 4688 11118 4968
rect 798 3608 11198 4688
rect 880 3328 11198 3608
rect 798 2143 11198 3328
<< metal4 >>
rect 2163 2128 2483 11472
rect 2823 2128 3143 11472
rect 4601 2128 4921 11472
rect 5261 2128 5581 11472
rect 7039 2128 7359 11472
rect 7699 2128 8019 11472
rect 9477 2128 9797 11472
rect 10137 2128 10457 11472
<< metal5 >>
rect 1056 10764 10904 11084
rect 1056 10104 10904 10424
rect 1056 8453 10904 8773
rect 1056 7793 10904 8113
rect 1056 6142 10904 6462
rect 1056 5482 10904 5802
rect 1056 3831 10904 4151
rect 1056 3171 10904 3491
<< labels >>
rlabel metal4 s 2823 2128 3143 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5261 2128 5581 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7699 2128 8019 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10137 2128 10457 11472 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3831 10904 4151 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6142 10904 6462 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8453 10904 8773 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 10764 10904 11084 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2163 2128 2483 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4601 2128 4921 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7039 2128 7359 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9477 2128 9797 11472 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3171 10904 3491 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5482 10904 5802 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7793 10904 8113 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 10104 10904 10424 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 8390 0 8446 800 6 a[0]
port 3 nsew signal input
rlabel metal3 s 11198 4768 11998 4888 6 a[1]
port 4 nsew signal input
rlabel metal3 s 11198 8848 11998 8968 6 a[2]
port 5 nsew signal input
rlabel metal2 s 7746 13342 7802 14142 6 a[3]
port 6 nsew signal input
rlabel metal2 s 4526 13342 4582 14142 6 a[4]
port 7 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 a[5]
port 8 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 a[6]
port 9 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 a[7]
port 10 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 b[0]
port 11 nsew signal input
rlabel metal3 s 11198 5448 11998 5568 6 b[1]
port 12 nsew signal input
rlabel metal3 s 11198 8168 11998 8288 6 b[2]
port 13 nsew signal input
rlabel metal2 s 7102 13342 7158 14142 6 b[3]
port 14 nsew signal input
rlabel metal2 s 3882 13342 3938 14142 6 b[4]
port 15 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 b[5]
port 16 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 b[6]
port 17 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 b[7]
port 18 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 cin
port 19 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 cout
port 20 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 op[0]
port 21 nsew signal input
rlabel metal3 s 11198 6808 11998 6928 6 op[1]
port 22 nsew signal input
rlabel metal3 s 11198 6128 11998 6248 6 op[2]
port 23 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 result[0]
port 24 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 result[1]
port 25 nsew signal output
rlabel metal3 s 11198 7488 11998 7608 6 result[2]
port 26 nsew signal output
rlabel metal2 s 5814 13342 5870 14142 6 result[3]
port 27 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 result[4]
port 28 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 result[5]
port 29 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 result[6]
port 30 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 result[7]
port 31 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 11998 14142
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 714904
string GDS_FILE /openlane/designs/alu_8bit/runs/RUN_2025.05.07_17.19.58/results/signoff/alu_8bit.magic.gds
string GDS_START 299672
<< end >>

