magic
tech sky130A
magscale 1 2
timestamp 1746638552
<< viali >>
rect 6561 11305 6595 11339
rect 8493 11237 8527 11271
rect 7113 11169 7147 11203
rect 4169 11101 4203 11135
rect 5365 11101 5399 11135
rect 5641 11101 5675 11135
rect 7389 11101 7423 11135
rect 8033 11101 8067 11135
rect 9137 11101 9171 11135
rect 6469 11033 6503 11067
rect 3985 10965 4019 10999
rect 4905 10965 4939 10999
rect 5457 10965 5491 10999
rect 8953 10965 8987 10999
rect 5073 10761 5107 10795
rect 5733 10761 5767 10795
rect 7297 10761 7331 10795
rect 8493 10761 8527 10795
rect 3985 10693 4019 10727
rect 5273 10693 5307 10727
rect 6193 10693 6227 10727
rect 1685 10625 1719 10659
rect 2053 10625 2087 10659
rect 2789 10625 2823 10659
rect 4169 10625 4203 10659
rect 4261 10625 4295 10659
rect 4537 10625 4571 10659
rect 4721 10625 4755 10659
rect 4813 10625 4847 10659
rect 5549 10625 5583 10659
rect 6009 10625 6043 10659
rect 6469 10625 6503 10659
rect 6653 10625 6687 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 8033 10625 8067 10659
rect 8677 10625 8711 10659
rect 2513 10557 2547 10591
rect 8217 10557 8251 10591
rect 1869 10489 1903 10523
rect 4905 10489 4939 10523
rect 1501 10421 1535 10455
rect 2605 10421 2639 10455
rect 2697 10421 2731 10455
rect 3985 10421 4019 10455
rect 4353 10421 4387 10455
rect 5089 10421 5123 10455
rect 5825 10421 5859 10455
rect 6561 10421 6595 10455
rect 6745 10421 6779 10455
rect 1501 10217 1535 10251
rect 4997 10217 5031 10251
rect 6009 10217 6043 10251
rect 5273 10149 5307 10183
rect 7573 10149 7607 10183
rect 2421 10081 2455 10115
rect 2881 10081 2915 10115
rect 3249 10081 3283 10115
rect 6653 10081 6687 10115
rect 1685 10013 1719 10047
rect 2145 10013 2179 10047
rect 2513 10013 2547 10047
rect 3433 10013 3467 10047
rect 3617 10013 3651 10047
rect 3893 10013 3927 10047
rect 3985 10013 4019 10047
rect 4353 10013 4387 10047
rect 4445 10013 4479 10047
rect 4629 10013 4663 10047
rect 4721 10013 4755 10047
rect 6193 10013 6227 10047
rect 6285 10013 6319 10047
rect 7113 10013 7147 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8033 10013 8067 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 1777 9945 1811 9979
rect 1869 9945 1903 9979
rect 2007 9945 2041 9979
rect 2789 9945 2823 9979
rect 5181 9945 5215 9979
rect 5457 9945 5491 9979
rect 6377 9945 6411 9979
rect 6495 9945 6529 9979
rect 6929 9945 6963 9979
rect 7941 9945 7975 9979
rect 8125 9945 8159 9979
rect 2237 9877 2271 9911
rect 4169 9877 4203 9911
rect 4813 9877 4847 9911
rect 4981 9877 5015 9911
rect 7297 9877 7331 9911
rect 2053 9673 2087 9707
rect 6377 9673 6411 9707
rect 2421 9605 2455 9639
rect 3801 9605 3835 9639
rect 7021 9605 7055 9639
rect 7297 9605 7331 9639
rect 2237 9537 2271 9571
rect 2973 9537 3007 9571
rect 3709 9537 3743 9571
rect 3893 9537 3927 9571
rect 4353 9537 4387 9571
rect 4905 9537 4939 9571
rect 6653 9537 6687 9571
rect 7573 9537 7607 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 8125 9537 8159 9571
rect 8309 9537 8343 9571
rect 2881 9469 2915 9503
rect 4721 9469 4755 9503
rect 4813 9469 4847 9503
rect 6561 9469 6595 9503
rect 6929 9469 6963 9503
rect 7205 9469 7239 9503
rect 7757 9469 7791 9503
rect 2605 9401 2639 9435
rect 8217 9401 8251 9435
rect 2789 9333 2823 9367
rect 7941 9333 7975 9367
rect 9873 9129 9907 9163
rect 9413 8993 9447 9027
rect 1409 8925 1443 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9505 8925 9539 8959
rect 10517 8925 10551 8959
rect 1593 8789 1627 8823
rect 10333 8789 10367 8823
rect 9689 8585 9723 8619
rect 9965 8517 9999 8551
rect 1685 8449 1719 8483
rect 2237 8449 2271 8483
rect 2421 8449 2455 8483
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 4721 8449 4755 8483
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 9413 8449 9447 8483
rect 10149 8449 10183 8483
rect 10241 8449 10275 8483
rect 4261 8381 4295 8415
rect 8953 8381 8987 8415
rect 9229 8381 9263 8415
rect 9321 8381 9355 8415
rect 9505 8381 9539 8415
rect 1501 8313 1535 8347
rect 2605 8313 2639 8347
rect 9781 8313 9815 8347
rect 10425 8313 10459 8347
rect 2053 8245 2087 8279
rect 4537 8245 4571 8279
rect 2973 8041 3007 8075
rect 3433 8041 3467 8075
rect 6561 8041 6595 8075
rect 6929 8041 6963 8075
rect 9597 8041 9631 8075
rect 10333 8041 10367 8075
rect 3249 7973 3283 8007
rect 2053 7905 2087 7939
rect 2329 7905 2363 7939
rect 2697 7905 2731 7939
rect 2789 7905 2823 7939
rect 4169 7905 4203 7939
rect 4629 7905 4663 7939
rect 4721 7905 4755 7939
rect 7757 7905 7791 7939
rect 8217 7905 8251 7939
rect 8309 7905 8343 7939
rect 1593 7837 1627 7871
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3801 7837 3835 7871
rect 5181 7837 5215 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 6009 7837 6043 7871
rect 6429 7837 6463 7871
rect 6745 7837 6779 7871
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 7389 7837 7423 7871
rect 7481 7837 7515 7871
rect 8033 7837 8067 7871
rect 8125 7837 8159 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 8953 7837 8987 7871
rect 9413 7837 9447 7871
rect 9689 7837 9723 7871
rect 10517 7837 10551 7871
rect 1685 7769 1719 7803
rect 1915 7769 1949 7803
rect 3401 7769 3435 7803
rect 3617 7769 3651 7803
rect 3893 7769 3927 7803
rect 6193 7769 6227 7803
rect 6285 7769 6319 7803
rect 9111 7769 9145 7803
rect 9229 7769 9263 7803
rect 9321 7769 9355 7803
rect 1409 7701 1443 7735
rect 2145 7701 2179 7735
rect 4353 7701 4387 7735
rect 4997 7701 5031 7735
rect 7849 7701 7883 7735
rect 8769 7701 8803 7735
rect 10149 7701 10183 7735
rect 1593 7497 1627 7531
rect 1777 7497 1811 7531
rect 2237 7497 2271 7531
rect 2789 7497 2823 7531
rect 4077 7497 4111 7531
rect 4445 7497 4479 7531
rect 6561 7497 6595 7531
rect 6745 7497 6779 7531
rect 7665 7497 7699 7531
rect 9045 7497 9079 7531
rect 2421 7429 2455 7463
rect 2605 7429 2639 7463
rect 3157 7429 3191 7463
rect 4537 7429 4571 7463
rect 4753 7429 4787 7463
rect 6193 7429 6227 7463
rect 8861 7429 8895 7463
rect 1409 7361 1443 7395
rect 1961 7361 1995 7395
rect 2973 7361 3007 7395
rect 3985 7361 4019 7395
rect 4261 7361 4295 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 6742 7361 6776 7395
rect 7113 7361 7147 7395
rect 7297 7361 7331 7395
rect 7757 7361 7791 7395
rect 8585 7361 8619 7395
rect 8769 7361 8803 7395
rect 9137 7361 9171 7395
rect 9413 7361 9447 7395
rect 9597 7361 9631 7395
rect 10425 7361 10459 7395
rect 7205 7293 7239 7327
rect 8677 7293 8711 7327
rect 9873 7293 9907 7327
rect 4905 7225 4939 7259
rect 7389 7225 7423 7259
rect 8861 7225 8895 7259
rect 9505 7225 9539 7259
rect 4721 7157 4755 7191
rect 8953 6953 8987 6987
rect 6469 6885 6503 6919
rect 9321 6817 9355 6851
rect 10333 6817 10367 6851
rect 5549 6749 5583 6783
rect 6009 6749 6043 6783
rect 6101 6749 6135 6783
rect 6745 6749 6779 6783
rect 6929 6749 6963 6783
rect 9137 6749 9171 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 7297 6681 7331 6715
rect 5917 6613 5951 6647
rect 6561 6613 6595 6647
rect 9689 6613 9723 6647
rect 4369 6409 4403 6443
rect 9045 6409 9079 6443
rect 2237 6341 2271 6375
rect 2421 6341 2455 6375
rect 4169 6341 4203 6375
rect 9873 6341 9907 6375
rect 1409 6273 1443 6307
rect 5365 6273 5399 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 9321 6273 9355 6307
rect 10425 6273 10459 6307
rect 5273 6205 5307 6239
rect 9137 6205 9171 6239
rect 9689 6205 9723 6239
rect 1593 6137 1627 6171
rect 9597 6137 9631 6171
rect 2053 6069 2087 6103
rect 4353 6069 4387 6103
rect 4537 6069 4571 6103
rect 4813 6069 4847 6103
rect 5457 6069 5491 6103
rect 9413 5865 9447 5899
rect 9965 5797 9999 5831
rect 10333 5797 10367 5831
rect 2053 5729 2087 5763
rect 2697 5729 2731 5763
rect 2789 5729 2823 5763
rect 2881 5729 2915 5763
rect 3065 5729 3099 5763
rect 4353 5729 4387 5763
rect 4721 5729 4755 5763
rect 4813 5729 4847 5763
rect 7941 5729 7975 5763
rect 10149 5729 10183 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 2421 5661 2455 5695
rect 3157 5661 3191 5695
rect 3433 5661 3467 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 4905 5661 4939 5695
rect 5181 5661 5215 5695
rect 5273 5661 5307 5695
rect 5457 5661 5491 5695
rect 5549 5661 5583 5695
rect 6745 5661 6779 5695
rect 6929 5661 6963 5695
rect 7205 5661 7239 5695
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 8309 5661 8343 5695
rect 8953 5661 8987 5695
rect 9597 5661 9631 5695
rect 9965 5661 9999 5695
rect 10517 5661 10551 5695
rect 1685 5593 1719 5627
rect 1777 5593 1811 5627
rect 1915 5593 1949 5627
rect 3249 5593 3283 5627
rect 4261 5593 4295 5627
rect 6837 5593 6871 5627
rect 7067 5593 7101 5627
rect 8125 5593 8159 5627
rect 8401 5593 8435 5627
rect 8585 5593 8619 5627
rect 1409 5525 1443 5559
rect 2145 5525 2179 5559
rect 2881 5525 2915 5559
rect 3617 5525 3651 5559
rect 3893 5525 3927 5559
rect 5733 5525 5767 5559
rect 6561 5525 6595 5559
rect 7757 5525 7791 5559
rect 8769 5525 8803 5559
rect 1501 5321 1535 5355
rect 2329 5321 2363 5355
rect 3617 5321 3651 5355
rect 4461 5321 4495 5355
rect 4629 5321 4663 5355
rect 6745 5321 6779 5355
rect 7481 5321 7515 5355
rect 10333 5321 10367 5355
rect 3801 5253 3835 5287
rect 4261 5253 4295 5287
rect 7849 5253 7883 5287
rect 1685 5185 1719 5219
rect 1961 5185 1995 5219
rect 2697 5185 2731 5219
rect 3525 5185 3559 5219
rect 3709 5185 3743 5219
rect 3985 5185 4019 5219
rect 4077 5185 4111 5219
rect 6469 5185 6503 5219
rect 7021 5185 7055 5219
rect 7297 5185 7331 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 9045 5185 9079 5219
rect 10517 5185 10551 5219
rect 2605 5117 2639 5151
rect 6929 5117 6963 5151
rect 7389 5117 7423 5151
rect 1777 5049 1811 5083
rect 3801 5049 3835 5083
rect 6653 5049 6687 5083
rect 9321 5049 9355 5083
rect 2697 4981 2731 5015
rect 4445 4981 4479 5015
rect 1593 4777 1627 4811
rect 6009 4777 6043 4811
rect 8033 4777 8067 4811
rect 9045 4709 9079 4743
rect 6653 4641 6687 4675
rect 7297 4641 7331 4675
rect 8217 4641 8251 4675
rect 8769 4641 8803 4675
rect 9505 4641 9539 4675
rect 1409 4573 1443 4607
rect 6101 4573 6135 4607
rect 6469 4573 6503 4607
rect 6929 4573 6963 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 8401 4573 8435 4607
rect 8677 4573 8711 4607
rect 7757 4437 7791 4471
rect 5517 4165 5551 4199
rect 5733 4165 5767 4199
rect 4261 4097 4295 4131
rect 4445 4097 4479 4131
rect 5825 4097 5859 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 8953 4097 8987 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 5273 4029 5307 4063
rect 7573 4029 7607 4063
rect 8217 4029 8251 4063
rect 8677 4029 8711 4063
rect 7113 3961 7147 3995
rect 4353 3893 4387 3927
rect 4813 3893 4847 3927
rect 5365 3893 5399 3927
rect 5549 3893 5583 3927
rect 5825 3893 5859 3927
rect 9597 3893 9631 3927
rect 4721 3689 4755 3723
rect 7481 3621 7515 3655
rect 7573 3621 7607 3655
rect 1501 3553 1535 3587
rect 2513 3553 2547 3587
rect 3157 3553 3191 3587
rect 3525 3553 3559 3587
rect 5457 3553 5491 3587
rect 5549 3553 5583 3587
rect 5917 3553 5951 3587
rect 6929 3553 6963 3587
rect 8769 3553 8803 3587
rect 10241 3553 10275 3587
rect 2053 3485 2087 3519
rect 2605 3485 2639 3519
rect 2697 3485 2731 3519
rect 2789 3485 2823 3519
rect 3249 3485 3283 3519
rect 4353 3485 4387 3519
rect 4445 3485 4479 3519
rect 4721 3485 4755 3519
rect 5825 3485 5859 3519
rect 6009 3485 6043 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 8585 3485 8619 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 9689 3485 9723 3519
rect 9882 3485 9916 3519
rect 3617 3417 3651 3451
rect 3985 3417 4019 3451
rect 4169 3417 4203 3451
rect 2329 3349 2363 3383
rect 2973 3349 3007 3383
rect 4997 3349 5031 3383
rect 5089 3349 5123 3383
rect 5733 3349 5767 3383
rect 7021 3349 7055 3383
rect 7113 3349 7147 3383
rect 7757 3349 7791 3383
rect 2053 3145 2087 3179
rect 2789 3145 2823 3179
rect 3985 3145 4019 3179
rect 4537 3145 4571 3179
rect 5457 3145 5491 3179
rect 7021 3145 7055 3179
rect 7849 3145 7883 3179
rect 8769 3145 8803 3179
rect 9137 3145 9171 3179
rect 9873 3145 9907 3179
rect 4689 3077 4723 3111
rect 4905 3077 4939 3111
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 4261 3009 4295 3043
rect 4997 3009 5031 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 7205 3009 7239 3043
rect 7573 3009 7607 3043
rect 7849 3009 7883 3043
rect 8033 3009 8067 3043
rect 8769 3009 8803 3043
rect 8953 3009 8987 3043
rect 9689 3009 9723 3043
rect 9781 3009 9815 3043
rect 10241 3009 10275 3043
rect 10425 3009 10459 3043
rect 3249 2941 3283 2975
rect 3985 2941 4019 2975
rect 7481 2941 7515 2975
rect 8401 2941 8435 2975
rect 9597 2941 9631 2975
rect 10149 2941 10183 2975
rect 10333 2941 10367 2975
rect 3157 2873 3191 2907
rect 7389 2873 7423 2907
rect 9321 2873 9355 2907
rect 4169 2805 4203 2839
rect 4721 2805 4755 2839
rect 7757 2805 7791 2839
rect 4169 2601 4203 2635
rect 4721 2601 4755 2635
rect 6745 2601 6779 2635
rect 8677 2601 8711 2635
rect 9321 2601 9355 2635
rect 9965 2601 9999 2635
rect 3985 2397 4019 2431
rect 4537 2397 4571 2431
rect 5457 2397 5491 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 8493 2397 8527 2431
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 5089 2329 5123 2363
rect 7389 2261 7423 2295
rect 8033 2261 8067 2295
<< metal1 >>
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 8202 11880 8208 11892
rect 7156 11852 8208 11880
rect 7156 11840 7162 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 1104 11450 10856 11472
rect 1104 11398 2169 11450
rect 2221 11398 2233 11450
rect 2285 11398 2297 11450
rect 2349 11398 2361 11450
rect 2413 11398 2425 11450
rect 2477 11398 4607 11450
rect 4659 11398 4671 11450
rect 4723 11398 4735 11450
rect 4787 11398 4799 11450
rect 4851 11398 4863 11450
rect 4915 11398 7045 11450
rect 7097 11398 7109 11450
rect 7161 11398 7173 11450
rect 7225 11398 7237 11450
rect 7289 11398 7301 11450
rect 7353 11398 9483 11450
rect 9535 11398 9547 11450
rect 9599 11398 9611 11450
rect 9663 11398 9675 11450
rect 9727 11398 9739 11450
rect 9791 11398 10856 11450
rect 1104 11376 10856 11398
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5868 11308 6561 11336
rect 5868 11296 5874 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 8481 11271 8539 11277
rect 8481 11268 8493 11271
rect 7116 11240 8493 11268
rect 7116 11212 7144 11240
rect 8481 11237 8493 11240
rect 8527 11237 8539 11271
rect 8481 11231 8539 11237
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 4580 11172 5672 11200
rect 4580 11160 4586 11172
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 3936 11104 4169 11132
rect 3936 11092 3942 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 5644 11141 5672 11172
rect 7098 11160 7104 11212
rect 7156 11160 7162 11212
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 5224 11104 5365 11132
rect 5224 11092 5230 11104
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7524 11104 8033 11132
rect 7524 11092 7530 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8260 11104 9137 11132
rect 8260 11092 8266 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 6454 11024 6460 11076
rect 6512 11024 6518 11076
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 3973 10999 4031 11005
rect 3973 10996 3985 10999
rect 3936 10968 3985 10996
rect 3936 10956 3942 10968
rect 3973 10965 3985 10968
rect 4019 10965 4031 10999
rect 3973 10959 4031 10965
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4893 10999 4951 11005
rect 4893 10996 4905 10999
rect 4304 10968 4905 10996
rect 4304 10956 4310 10968
rect 4893 10965 4905 10968
rect 4939 10965 4951 10999
rect 4893 10959 4951 10965
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 5132 10968 5457 10996
rect 5132 10956 5138 10968
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5445 10959 5503 10965
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8941 10999 8999 11005
rect 8941 10996 8953 10999
rect 8352 10968 8953 10996
rect 8352 10956 8358 10968
rect 8941 10965 8953 10968
rect 8987 10965 8999 10999
rect 8941 10959 8999 10965
rect 1104 10906 10856 10928
rect 1104 10854 2829 10906
rect 2881 10854 2893 10906
rect 2945 10854 2957 10906
rect 3009 10854 3021 10906
rect 3073 10854 3085 10906
rect 3137 10854 5267 10906
rect 5319 10854 5331 10906
rect 5383 10854 5395 10906
rect 5447 10854 5459 10906
rect 5511 10854 5523 10906
rect 5575 10854 7705 10906
rect 7757 10854 7769 10906
rect 7821 10854 7833 10906
rect 7885 10854 7897 10906
rect 7949 10854 7961 10906
rect 8013 10854 10143 10906
rect 10195 10854 10207 10906
rect 10259 10854 10271 10906
rect 10323 10854 10335 10906
rect 10387 10854 10399 10906
rect 10451 10854 10856 10906
rect 1104 10832 10856 10854
rect 5074 10801 5080 10804
rect 5061 10795 5080 10801
rect 5061 10792 5073 10795
rect 4632 10764 5073 10792
rect 3418 10684 3424 10736
rect 3476 10724 3482 10736
rect 3973 10727 4031 10733
rect 3973 10724 3985 10727
rect 3476 10696 3985 10724
rect 3476 10684 3482 10696
rect 3973 10693 3985 10696
rect 4019 10724 4031 10727
rect 4632 10724 4660 10764
rect 5061 10761 5073 10764
rect 5061 10755 5080 10761
rect 5074 10752 5080 10755
rect 5132 10752 5138 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 6454 10792 6460 10804
rect 5767 10764 6460 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 7098 10792 7104 10804
rect 6564 10764 7104 10792
rect 4019 10696 4660 10724
rect 4019 10693 4031 10696
rect 3973 10687 4031 10693
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1719 10628 1900 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1872 10529 1900 10628
rect 2038 10616 2044 10668
rect 2096 10616 2102 10668
rect 2774 10616 2780 10668
rect 2832 10616 2838 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3878 10588 3884 10600
rect 2547 10560 3884 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4172 10588 4200 10619
rect 4246 10616 4252 10668
rect 4304 10616 4310 10668
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 4632 10656 4660 10696
rect 5258 10684 5264 10736
rect 5316 10684 5322 10736
rect 6181 10727 6239 10733
rect 6181 10693 6193 10727
rect 6227 10724 6239 10727
rect 6564 10724 6592 10764
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7285 10795 7343 10801
rect 7285 10761 7297 10795
rect 7331 10792 7343 10795
rect 7466 10792 7472 10804
rect 7331 10764 7472 10792
rect 7331 10761 7343 10764
rect 7285 10755 7343 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10761 8539 10795
rect 8481 10755 8539 10761
rect 7374 10724 7380 10736
rect 6227 10696 6592 10724
rect 6656 10696 7380 10724
rect 6227 10693 6239 10696
rect 6181 10687 6239 10693
rect 4571 10628 4660 10656
rect 4709 10659 4767 10665
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 5276 10656 5304 10684
rect 4847 10628 5304 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 4724 10588 4752 10619
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 6656 10665 6684 10696
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 8202 10724 8208 10736
rect 8036 10696 8208 10724
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 6457 10659 6515 10665
rect 6457 10656 6469 10659
rect 6043 10628 6469 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6457 10625 6469 10628
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 4172 10560 5120 10588
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10489 1915 10523
rect 1857 10483 1915 10489
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 4893 10523 4951 10529
rect 4893 10520 4905 10523
rect 4120 10492 4905 10520
rect 4120 10480 4126 10492
rect 4893 10489 4905 10492
rect 4939 10489 4951 10523
rect 4893 10483 4951 10489
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 900 10424 1501 10452
rect 900 10412 906 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 1728 10424 2605 10452
rect 1728 10412 1734 10424
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 2593 10415 2651 10421
rect 2685 10455 2743 10461
rect 2685 10421 2697 10455
rect 2731 10452 2743 10455
rect 3234 10452 3240 10464
rect 2731 10424 3240 10452
rect 2731 10421 2743 10424
rect 2685 10415 2743 10421
rect 3234 10412 3240 10424
rect 3292 10452 3298 10464
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3292 10424 3985 10452
rect 3292 10412 3298 10424
rect 3973 10421 3985 10424
rect 4019 10421 4031 10455
rect 3973 10415 4031 10421
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4430 10452 4436 10464
rect 4387 10424 4436 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 5092 10461 5120 10560
rect 6472 10520 6500 10619
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7116 10588 7144 10619
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 8036 10665 8064 10696
rect 8202 10684 8208 10696
rect 8260 10724 8266 10736
rect 8496 10724 8524 10755
rect 8260 10696 8524 10724
rect 8260 10684 8266 10696
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7708 10628 8033 10656
rect 7708 10616 7714 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8168 10628 8677 10656
rect 8168 10616 8174 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 7374 10588 7380 10600
rect 7116 10560 7380 10588
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 8570 10588 8576 10600
rect 8251 10560 8576 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8294 10520 8300 10532
rect 6472 10492 8300 10520
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5350 10452 5356 10464
rect 5123 10424 5356 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5810 10412 5816 10464
rect 5868 10412 5874 10464
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6236 10424 6561 10452
rect 6236 10412 6242 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 6733 10455 6791 10461
rect 6733 10452 6745 10455
rect 6696 10424 6745 10452
rect 6696 10412 6702 10424
rect 6733 10421 6745 10424
rect 6779 10421 6791 10455
rect 6733 10415 6791 10421
rect 1104 10362 10856 10384
rect 1104 10310 2169 10362
rect 2221 10310 2233 10362
rect 2285 10310 2297 10362
rect 2349 10310 2361 10362
rect 2413 10310 2425 10362
rect 2477 10310 4607 10362
rect 4659 10310 4671 10362
rect 4723 10310 4735 10362
rect 4787 10310 4799 10362
rect 4851 10310 4863 10362
rect 4915 10310 7045 10362
rect 7097 10310 7109 10362
rect 7161 10310 7173 10362
rect 7225 10310 7237 10362
rect 7289 10310 7301 10362
rect 7353 10310 9483 10362
rect 9535 10310 9547 10362
rect 9599 10310 9611 10362
rect 9663 10310 9675 10362
rect 9727 10310 9739 10362
rect 9791 10310 10856 10362
rect 1104 10288 10856 10310
rect 1489 10251 1547 10257
rect 1489 10217 1501 10251
rect 1535 10248 1547 10251
rect 2038 10248 2044 10260
rect 1535 10220 2044 10248
rect 1535 10217 1547 10220
rect 1489 10211 1547 10217
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 4985 10251 5043 10257
rect 4985 10248 4997 10251
rect 3844 10220 4997 10248
rect 3844 10208 3850 10220
rect 4985 10217 4997 10220
rect 5031 10217 5043 10251
rect 4985 10211 5043 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5592 10220 6009 10248
rect 5592 10208 5598 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 6328 10220 8064 10248
rect 6328 10208 6334 10220
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 4062 10180 4068 10192
rect 2832 10152 4068 10180
rect 2832 10140 2838 10152
rect 4062 10140 4068 10152
rect 4120 10180 4126 10192
rect 4120 10152 4660 10180
rect 4120 10140 4126 10152
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 1452 10084 2421 10112
rect 1452 10072 1458 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 2409 10075 2467 10081
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3237 10115 3295 10121
rect 3237 10112 3249 10115
rect 2915 10084 3249 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3237 10081 3249 10084
rect 3283 10112 3295 10115
rect 4154 10112 4160 10124
rect 3283 10084 4160 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 4632 10112 4660 10152
rect 5258 10140 5264 10192
rect 5316 10140 5322 10192
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 7561 10183 7619 10189
rect 7561 10180 7573 10183
rect 5408 10152 7573 10180
rect 5408 10140 5414 10152
rect 7561 10149 7573 10152
rect 7607 10149 7619 10183
rect 7561 10143 7619 10149
rect 5368 10112 5396 10140
rect 4632 10084 4752 10112
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 2130 10004 2136 10056
rect 2188 10004 2194 10056
rect 2498 10004 2504 10056
rect 2556 10004 2562 10056
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10044 3663 10047
rect 3878 10044 3884 10056
rect 3651 10016 3884 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 4019 10016 4353 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 4341 10013 4353 10016
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4724 10053 4752 10084
rect 5276 10084 5396 10112
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 1762 9936 1768 9988
rect 1820 9936 1826 9988
rect 1854 9936 1860 9988
rect 1912 9936 1918 9988
rect 1995 9979 2053 9985
rect 1995 9945 2007 9979
rect 2041 9976 2053 9979
rect 2777 9979 2835 9985
rect 2041 9948 2268 9976
rect 2041 9945 2053 9948
rect 1995 9939 2053 9945
rect 2240 9917 2268 9948
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 3326 9976 3332 9988
rect 2823 9948 3332 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3326 9936 3332 9948
rect 3384 9936 3390 9988
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5276 9976 5304 10084
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 5868 10084 6316 10112
rect 5868 10072 5874 10084
rect 6178 10004 6184 10056
rect 6236 10004 6242 10056
rect 6288 10053 6316 10084
rect 6638 10072 6644 10124
rect 6696 10072 6702 10124
rect 7650 10112 7656 10124
rect 7116 10084 7656 10112
rect 7116 10053 7144 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 8036 10053 8064 10220
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7524 10016 7573 10044
rect 7524 10004 7530 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8021 10047 8079 10053
rect 7791 10016 7880 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 5215 9948 5304 9976
rect 5445 9979 5503 9985
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 5445 9945 5457 9979
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9877 2283 9911
rect 2225 9871 2283 9877
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9908 4215 9911
rect 4246 9908 4252 9920
rect 4203 9880 4252 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 4798 9868 4804 9920
rect 4856 9868 4862 9920
rect 4969 9911 5027 9917
rect 4969 9877 4981 9911
rect 5015 9908 5027 9911
rect 5460 9908 5488 9939
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 6365 9979 6423 9985
rect 6365 9976 6377 9979
rect 5960 9948 6377 9976
rect 5960 9936 5966 9948
rect 6365 9945 6377 9948
rect 6411 9945 6423 9979
rect 6365 9939 6423 9945
rect 6454 9936 6460 9988
rect 6512 9985 6518 9988
rect 6512 9979 6541 9985
rect 6529 9945 6541 9979
rect 6512 9939 6541 9945
rect 6917 9979 6975 9985
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 7852 9976 7880 10016
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8260 10016 8401 10044
rect 8260 10004 8266 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 6963 9948 7880 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 6512 9936 6518 9939
rect 6822 9908 6828 9920
rect 5015 9880 6828 9908
rect 5015 9877 5027 9880
rect 4969 9871 5027 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 7064 9880 7297 9908
rect 7064 9868 7070 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7852 9908 7880 9948
rect 7929 9979 7987 9985
rect 7929 9945 7941 9979
rect 7975 9976 7987 9979
rect 8113 9979 8171 9985
rect 8113 9976 8125 9979
rect 7975 9948 8125 9976
rect 7975 9945 7987 9948
rect 7929 9939 7987 9945
rect 8113 9945 8125 9948
rect 8159 9945 8171 9979
rect 8113 9939 8171 9945
rect 8294 9908 8300 9920
rect 7852 9880 8300 9908
rect 7285 9871 7343 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 1104 9818 10856 9840
rect 1104 9766 2829 9818
rect 2881 9766 2893 9818
rect 2945 9766 2957 9818
rect 3009 9766 3021 9818
rect 3073 9766 3085 9818
rect 3137 9766 5267 9818
rect 5319 9766 5331 9818
rect 5383 9766 5395 9818
rect 5447 9766 5459 9818
rect 5511 9766 5523 9818
rect 5575 9766 7705 9818
rect 7757 9766 7769 9818
rect 7821 9766 7833 9818
rect 7885 9766 7897 9818
rect 7949 9766 7961 9818
rect 8013 9766 10143 9818
rect 10195 9766 10207 9818
rect 10259 9766 10271 9818
rect 10323 9766 10335 9818
rect 10387 9766 10399 9818
rect 10451 9766 10856 9818
rect 1104 9744 10856 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 2130 9704 2136 9716
rect 2087 9676 2136 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 5626 9704 5632 9716
rect 4672 9676 5632 9704
rect 4672 9664 4678 9676
rect 5626 9664 5632 9676
rect 5684 9704 5690 9716
rect 6270 9704 6276 9716
rect 5684 9676 6276 9704
rect 5684 9664 5690 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6365 9707 6423 9713
rect 6365 9673 6377 9707
rect 6411 9704 6423 9707
rect 6454 9704 6460 9716
rect 6411 9676 6460 9704
rect 6411 9673 6423 9676
rect 6365 9667 6423 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 7024 9676 8064 9704
rect 7024 9648 7052 9676
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2498 9636 2504 9648
rect 2455 9608 2504 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 2498 9596 2504 9608
rect 2556 9636 2562 9648
rect 3786 9636 3792 9648
rect 2556 9608 3792 9636
rect 2556 9596 2562 9608
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 4798 9596 4804 9648
rect 4856 9596 4862 9648
rect 7006 9596 7012 9648
rect 7064 9596 7070 9648
rect 7285 9639 7343 9645
rect 7285 9605 7297 9639
rect 7331 9636 7343 9639
rect 7331 9608 7880 9636
rect 7331 9605 7343 9608
rect 7285 9599 7343 9605
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 2004 9540 2237 9568
rect 2004 9528 2010 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3234 9568 3240 9580
rect 3007 9540 3240 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3476 9540 3709 9568
rect 3476 9528 3482 9540
rect 3697 9537 3709 9540
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3878 9528 3884 9580
rect 3936 9528 3942 9580
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4341 9571 4399 9577
rect 4341 9568 4353 9571
rect 4212 9540 4353 9568
rect 4212 9528 4218 9540
rect 4341 9537 4353 9540
rect 4387 9537 4399 9571
rect 4816 9568 4844 9596
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4816 9540 4905 9568
rect 4341 9531 4399 9537
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7374 9568 7380 9580
rect 6687 9540 7380 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7374 9528 7380 9540
rect 7432 9568 7438 9580
rect 7852 9577 7880 9608
rect 8036 9577 8064 9676
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7432 9540 7573 9568
rect 7432 9528 7438 9540
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8202 9568 8208 9580
rect 8159 9540 8208 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9500 2927 9503
rect 3896 9500 3924 9528
rect 2915 9472 3924 9500
rect 4709 9503 4767 9509
rect 2915 9469 2927 9472
rect 2869 9463 2927 9469
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9500 4859 9503
rect 5074 9500 5080 9512
rect 4847 9472 5080 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 1762 9392 1768 9444
rect 1820 9432 1826 9444
rect 2593 9435 2651 9441
rect 2593 9432 2605 9435
rect 1820 9404 2605 9432
rect 1820 9392 1826 9404
rect 2593 9401 2605 9404
rect 2639 9401 2651 9435
rect 4724 9432 4752 9463
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6512 9472 6561 9500
rect 6512 9460 6518 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6880 9472 6929 9500
rect 6880 9460 6886 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 4982 9432 4988 9444
rect 4724 9404 4988 9432
rect 2593 9395 2651 9401
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 5092 9432 5120 9460
rect 7208 9432 7236 9463
rect 5092 9404 7236 9432
rect 7576 9432 7604 9531
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 8570 9500 8576 9512
rect 7791 9472 8576 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7576 9404 8217 9432
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 2774 9324 2780 9376
rect 2832 9324 2838 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 6822 9364 6828 9376
rect 3384 9336 6828 9364
rect 3384 9324 3390 9336
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 6972 9336 7941 9364
rect 6972 9324 6978 9336
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 7929 9327 7987 9333
rect 1104 9274 10856 9296
rect 1104 9222 2169 9274
rect 2221 9222 2233 9274
rect 2285 9222 2297 9274
rect 2349 9222 2361 9274
rect 2413 9222 2425 9274
rect 2477 9222 4607 9274
rect 4659 9222 4671 9274
rect 4723 9222 4735 9274
rect 4787 9222 4799 9274
rect 4851 9222 4863 9274
rect 4915 9222 7045 9274
rect 7097 9222 7109 9274
rect 7161 9222 7173 9274
rect 7225 9222 7237 9274
rect 7289 9222 7301 9274
rect 7353 9222 9483 9274
rect 9535 9222 9547 9274
rect 9599 9222 9611 9274
rect 9663 9222 9675 9274
rect 9727 9222 9739 9274
rect 9791 9222 10856 9274
rect 1104 9200 10856 9222
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 8628 9132 9873 9160
rect 8628 9120 8634 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 9861 9123 9919 9129
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 5684 8996 9413 9024
rect 5684 8984 5690 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 9508 8888 9536 8919
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 9456 8860 9536 8888
rect 9456 8848 9462 8860
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 3234 8820 3240 8832
rect 1627 8792 3240 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9858 8820 9864 8832
rect 9088 8792 9864 8820
rect 9088 8780 9094 8792
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10321 8823 10379 8829
rect 10321 8820 10333 8823
rect 10008 8792 10333 8820
rect 10008 8780 10014 8792
rect 10321 8789 10333 8792
rect 10367 8789 10379 8823
rect 10321 8783 10379 8789
rect 1104 8730 10856 8752
rect 1104 8678 2829 8730
rect 2881 8678 2893 8730
rect 2945 8678 2957 8730
rect 3009 8678 3021 8730
rect 3073 8678 3085 8730
rect 3137 8678 5267 8730
rect 5319 8678 5331 8730
rect 5383 8678 5395 8730
rect 5447 8678 5459 8730
rect 5511 8678 5523 8730
rect 5575 8678 7705 8730
rect 7757 8678 7769 8730
rect 7821 8678 7833 8730
rect 7885 8678 7897 8730
rect 7949 8678 7961 8730
rect 8013 8678 10143 8730
rect 10195 8678 10207 8730
rect 10259 8678 10271 8730
rect 10323 8678 10335 8730
rect 10387 8678 10399 8730
rect 10451 8678 10856 8730
rect 1104 8656 10856 8678
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 9180 8588 9689 8616
rect 9180 8576 9186 8588
rect 9677 8585 9689 8588
rect 9723 8585 9735 8619
rect 9677 8579 9735 8585
rect 9950 8548 9956 8560
rect 8864 8520 9956 8548
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 2004 8452 2237 8480
rect 2004 8440 2010 8452
rect 2225 8449 2237 8452
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2406 8440 2412 8492
rect 2464 8440 2470 8492
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2516 8412 2544 8443
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2648 8452 2697 8480
rect 2648 8440 2654 8452
rect 2685 8449 2697 8452
rect 2731 8480 2743 8483
rect 4709 8483 4767 8489
rect 2731 8452 4292 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 4264 8421 4292 8452
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 5166 8480 5172 8492
rect 4755 8452 5172 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8864 8489 8892 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8720 8452 8861 8480
rect 8720 8440 8726 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9582 8480 9588 8492
rect 9447 8452 9588 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9916 8452 10149 8480
rect 9916 8440 9922 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 4249 8415 4307 8421
rect 2516 8384 2728 8412
rect 2700 8356 2728 8384
rect 4249 8381 4261 8415
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 8987 8384 9229 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9306 8372 9312 8424
rect 9364 8372 9370 8424
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 1636 8316 2605 8344
rect 1636 8304 1642 8316
rect 2593 8313 2605 8316
rect 2639 8313 2651 8347
rect 2593 8307 2651 8313
rect 2682 8304 2688 8356
rect 2740 8304 2746 8356
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 9769 8347 9827 8353
rect 9769 8344 9781 8347
rect 8628 8316 9781 8344
rect 8628 8304 8634 8316
rect 9769 8313 9781 8316
rect 9815 8313 9827 8347
rect 9769 8307 9827 8313
rect 10413 8347 10471 8353
rect 10413 8313 10425 8347
rect 10459 8344 10471 8347
rect 10686 8344 10692 8356
rect 10459 8316 10692 8344
rect 10459 8313 10471 8316
rect 10413 8307 10471 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 2038 8236 2044 8288
rect 2096 8236 2102 8288
rect 4522 8236 4528 8288
rect 4580 8236 4586 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9490 8276 9496 8288
rect 9088 8248 9496 8276
rect 9088 8236 9094 8248
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 9950 8276 9956 8288
rect 9640 8248 9956 8276
rect 9640 8236 9646 8248
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 1104 8186 10856 8208
rect 1104 8134 2169 8186
rect 2221 8134 2233 8186
rect 2285 8134 2297 8186
rect 2349 8134 2361 8186
rect 2413 8134 2425 8186
rect 2477 8134 4607 8186
rect 4659 8134 4671 8186
rect 4723 8134 4735 8186
rect 4787 8134 4799 8186
rect 4851 8134 4863 8186
rect 4915 8134 7045 8186
rect 7097 8134 7109 8186
rect 7161 8134 7173 8186
rect 7225 8134 7237 8186
rect 7289 8134 7301 8186
rect 7353 8134 9483 8186
rect 9535 8134 9547 8186
rect 9599 8134 9611 8186
rect 9663 8134 9675 8186
rect 9727 8134 9739 8186
rect 9791 8134 10856 8186
rect 1104 8112 10856 8134
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2958 8072 2964 8084
rect 2556 8044 2964 8072
rect 2556 8032 2562 8044
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3326 8072 3332 8084
rect 3068 8044 3332 8072
rect 1394 7964 1400 8016
rect 1452 8004 1458 8016
rect 2130 8004 2136 8016
rect 1452 7976 2136 8004
rect 1452 7964 1458 7976
rect 2130 7964 2136 7976
rect 2188 8004 2194 8016
rect 3068 8004 3096 8044
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 4246 8072 4252 8084
rect 3467 8044 4252 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6822 8072 6828 8084
rect 6595 8044 6828 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 6963 8044 9168 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 2188 7976 2360 8004
rect 2188 7964 2194 7976
rect 1854 7936 1860 7948
rect 1780 7908 1860 7936
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 1780 7877 1808 7908
rect 1854 7896 1860 7908
rect 1912 7896 1918 7948
rect 2038 7896 2044 7948
rect 2096 7896 2102 7948
rect 2332 7945 2360 7976
rect 2700 7976 3096 8004
rect 3237 8007 3295 8013
rect 2700 7945 2728 7976
rect 3237 7973 3249 8007
rect 3283 8004 3295 8007
rect 3283 7976 4752 8004
rect 3283 7973 3295 7976
rect 3237 7967 3295 7973
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7905 2375 7939
rect 2317 7899 2375 7905
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7905 2743 7939
rect 2685 7899 2743 7905
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 4157 7939 4215 7945
rect 4157 7936 4169 7939
rect 2823 7908 4169 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 3252 7880 3280 7908
rect 4157 7905 4169 7908
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 4614 7896 4620 7948
rect 4672 7896 4678 7948
rect 4724 7945 4752 7976
rect 6454 7964 6460 8016
rect 6512 7964 6518 8016
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 8018 8004 8024 8016
rect 6788 7976 8024 8004
rect 6788 7964 6794 7976
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 9030 8004 9036 8016
rect 8128 7976 8340 8004
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 6472 7936 6500 7964
rect 7745 7939 7803 7945
rect 4709 7899 4767 7905
rect 5092 7908 5488 7936
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2498 7868 2504 7880
rect 2455 7840 2504 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2866 7828 2872 7880
rect 2924 7828 2930 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3142 7868 3148 7880
rect 3099 7840 3148 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3234 7828 3240 7880
rect 3292 7828 3298 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 5092 7868 5120 7908
rect 4580 7840 5120 7868
rect 4580 7828 4586 7840
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5460 7877 5488 7908
rect 6012 7908 7512 7936
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 5626 7868 5632 7880
rect 5583 7840 5632 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7769 1731 7803
rect 1673 7763 1731 7769
rect 1903 7803 1961 7809
rect 1903 7769 1915 7803
rect 1949 7800 1961 7803
rect 1949 7772 2176 7800
rect 1949 7769 1961 7772
rect 1903 7763 1961 7769
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 1578 7732 1584 7744
rect 1443 7704 1584 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 1688 7732 1716 7763
rect 2038 7732 2044 7744
rect 1688 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2148 7741 2176 7772
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 3389 7803 3447 7809
rect 3389 7800 3401 7803
rect 3016 7772 3401 7800
rect 3016 7760 3022 7772
rect 3389 7769 3401 7772
rect 3435 7769 3447 7803
rect 3389 7763 3447 7769
rect 3602 7760 3608 7812
rect 3660 7760 3666 7812
rect 3881 7803 3939 7809
rect 3881 7769 3893 7803
rect 3927 7800 3939 7803
rect 5276 7800 5304 7831
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 6012 7877 6040 7908
rect 6454 7877 6460 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5868 7840 6009 7868
rect 5868 7828 5874 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 5997 7831 6055 7837
rect 6417 7871 6460 7877
rect 6417 7837 6429 7871
rect 6417 7831 6460 7837
rect 6454 7828 6460 7831
rect 6512 7828 6518 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6604 7840 6745 7868
rect 6604 7828 6610 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 3927 7772 5304 7800
rect 3927 7769 3939 7772
rect 3881 7763 3939 7769
rect 6178 7760 6184 7812
rect 6236 7760 6242 7812
rect 6273 7803 6331 7809
rect 6273 7769 6285 7803
rect 6319 7800 6331 7803
rect 7300 7800 7328 7831
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 7484 7877 7512 7908
rect 7745 7905 7757 7939
rect 7791 7936 7803 7939
rect 8128 7936 8156 7976
rect 7791 7908 8156 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 8202 7896 8208 7948
rect 8260 7896 8266 7948
rect 8312 7945 8340 7976
rect 8772 7976 9036 8004
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7905 8355 7939
rect 8772 7936 8800 7976
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9140 8004 9168 8044
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 9456 8044 9597 8072
rect 9456 8032 9462 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 9916 8044 10333 8072
rect 9916 8032 9922 8044
rect 10321 8041 10333 8044
rect 10367 8041 10379 8075
rect 10321 8035 10379 8041
rect 10226 8004 10232 8016
rect 9140 7976 10232 8004
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 8297 7899 8355 7905
rect 8496 7908 8800 7936
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8386 7868 8392 7880
rect 8159 7840 8392 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8036 7800 8064 7831
rect 8386 7828 8392 7840
rect 8444 7868 8450 7880
rect 8496 7868 8524 7908
rect 8444 7840 8524 7868
rect 8444 7828 8450 7840
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 8772 7877 8800 7908
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 8904 7908 9076 7936
rect 8904 7896 8910 7908
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 9048 7868 9076 7908
rect 9401 7871 9459 7877
rect 9401 7870 9413 7871
rect 9324 7868 9413 7870
rect 9048 7842 9413 7868
rect 9048 7840 9352 7842
rect 8941 7831 8999 7837
rect 9401 7837 9413 7842
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 8588 7800 8616 7828
rect 6319 7772 6776 7800
rect 7300 7772 8616 7800
rect 6319 7769 6331 7772
rect 6273 7763 6331 7769
rect 6748 7744 6776 7772
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 8956 7800 8984 7831
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9548 7840 9689 7868
rect 9548 7828 9554 7840
rect 9677 7837 9689 7840
rect 9723 7868 9735 7871
rect 9950 7868 9956 7880
rect 9723 7840 9956 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 8720 7772 8984 7800
rect 9099 7803 9157 7809
rect 8720 7760 8726 7772
rect 9099 7769 9111 7803
rect 9145 7800 9157 7803
rect 9145 7769 9168 7800
rect 9099 7763 9168 7769
rect 2133 7735 2191 7741
rect 2133 7701 2145 7735
rect 2179 7701 2191 7735
rect 2133 7695 2191 7701
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4341 7735 4399 7741
rect 4341 7732 4353 7735
rect 4212 7704 4353 7732
rect 4212 7692 4218 7704
rect 4341 7701 4353 7704
rect 4387 7701 4399 7735
rect 4341 7695 4399 7701
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4488 7704 4997 7732
rect 4488 7692 4494 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 4985 7695 5043 7701
rect 6730 7692 6736 7744
rect 6788 7692 6794 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7156 7704 7849 7732
rect 7156 7692 7162 7704
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 8757 7735 8815 7741
rect 8757 7701 8769 7735
rect 8803 7732 8815 7735
rect 8846 7732 8852 7744
rect 8803 7704 8852 7732
rect 8803 7701 8815 7704
rect 8757 7695 8815 7701
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 9140 7732 9168 7763
rect 9214 7760 9220 7812
rect 9272 7760 9278 7812
rect 9306 7760 9312 7812
rect 9364 7760 9370 7812
rect 10042 7800 10048 7812
rect 9416 7772 10048 7800
rect 9416 7732 9444 7772
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 9140 7704 9444 7732
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 9548 7704 10149 7732
rect 9548 7692 9554 7704
rect 10137 7701 10149 7704
rect 10183 7701 10195 7735
rect 10137 7695 10195 7701
rect 1104 7642 10856 7664
rect 1104 7590 2829 7642
rect 2881 7590 2893 7642
rect 2945 7590 2957 7642
rect 3009 7590 3021 7642
rect 3073 7590 3085 7642
rect 3137 7590 5267 7642
rect 5319 7590 5331 7642
rect 5383 7590 5395 7642
rect 5447 7590 5459 7642
rect 5511 7590 5523 7642
rect 5575 7590 7705 7642
rect 7757 7590 7769 7642
rect 7821 7590 7833 7642
rect 7885 7590 7897 7642
rect 7949 7590 7961 7642
rect 8013 7590 10143 7642
rect 10195 7590 10207 7642
rect 10259 7590 10271 7642
rect 10323 7590 10335 7642
rect 10387 7590 10399 7642
rect 10451 7590 10856 7642
rect 1104 7568 10856 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 1596 7460 1624 7491
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 1765 7531 1823 7537
rect 1765 7528 1777 7531
rect 1728 7500 1777 7528
rect 1728 7488 1734 7500
rect 1765 7497 1777 7500
rect 1811 7497 1823 7531
rect 1765 7491 1823 7497
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 2096 7500 2237 7528
rect 2096 7488 2102 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 3234 7528 3240 7540
rect 2823 7500 3240 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 4065 7531 4123 7537
rect 3384 7500 4016 7528
rect 3384 7488 3390 7500
rect 2409 7463 2467 7469
rect 2409 7460 2421 7463
rect 1596 7432 2421 7460
rect 2409 7429 2421 7432
rect 2455 7429 2467 7463
rect 2409 7423 2467 7429
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 900 7364 1409 7392
rect 900 7352 906 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1636 7364 1961 7392
rect 1636 7352 1642 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 2424 7392 2452 7423
rect 2590 7420 2596 7472
rect 2648 7420 2654 7472
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 3145 7463 3203 7469
rect 3145 7460 3157 7463
rect 2740 7432 3157 7460
rect 2740 7420 2746 7432
rect 3145 7429 3157 7432
rect 3191 7460 3203 7463
rect 3786 7460 3792 7472
rect 3191 7432 3792 7460
rect 3191 7429 3203 7432
rect 3145 7423 3203 7429
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 3988 7460 4016 7500
rect 4065 7497 4077 7531
rect 4111 7528 4123 7531
rect 4246 7528 4252 7540
rect 4111 7500 4252 7528
rect 4111 7497 4123 7500
rect 4065 7491 4123 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 5166 7528 5172 7540
rect 4479 7500 5172 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 6733 7531 6791 7537
rect 6733 7497 6745 7531
rect 6779 7497 6791 7531
rect 6733 7491 6791 7497
rect 4525 7463 4583 7469
rect 4525 7460 4537 7463
rect 3988 7432 4537 7460
rect 2700 7392 2728 7420
rect 2424 7364 2728 7392
rect 2961 7395 3019 7401
rect 1949 7355 2007 7361
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3326 7392 3332 7404
rect 3007 7364 3332 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 4264 7401 4292 7432
rect 4525 7429 4537 7432
rect 4571 7429 4583 7463
rect 4741 7463 4799 7469
rect 4741 7460 4753 7463
rect 4525 7423 4583 7429
rect 4632 7432 4753 7460
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3660 7364 3985 7392
rect 3660 7352 3666 7364
rect 3973 7361 3985 7364
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 3988 7324 4016 7355
rect 4632 7324 4660 7432
rect 4741 7429 4753 7432
rect 4787 7460 4799 7463
rect 4982 7460 4988 7472
rect 4787 7432 4988 7460
rect 4787 7429 4799 7432
rect 4741 7423 4799 7429
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 6181 7463 6239 7469
rect 6181 7429 6193 7463
rect 6227 7460 6239 7463
rect 6748 7460 6776 7491
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7432 7500 7665 7528
rect 7432 7488 7438 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 9033 7531 9091 7537
rect 8720 7500 8984 7528
rect 8720 7488 8726 7500
rect 6227 7432 7328 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 5810 7352 5816 7404
rect 5868 7352 5874 7404
rect 5994 7352 6000 7404
rect 6052 7352 6058 7404
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7300 7401 7328 7432
rect 8846 7420 8852 7472
rect 8904 7420 8910 7472
rect 8956 7460 8984 7500
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9490 7528 9496 7540
rect 9079 7500 9496 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 8956 7432 9444 7460
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 8386 7392 8392 7404
rect 7791 7364 8392 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8570 7352 8576 7404
rect 8628 7352 8634 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 3988 7296 4660 7324
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 7006 7324 7012 7336
rect 6236 7296 7012 7324
rect 6236 7284 6242 7296
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 7239 7296 8677 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8772 7324 8800 7355
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 9088 7364 9137 7392
rect 9088 7352 9094 7364
rect 9125 7361 9137 7364
rect 9171 7392 9183 7395
rect 9214 7392 9220 7404
rect 9171 7364 9220 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9416 7401 9444 7432
rect 9858 7420 9864 7472
rect 9916 7420 9922 7472
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7392 9643 7395
rect 9876 7392 9904 7420
rect 10226 7392 10232 7404
rect 9631 7364 10232 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 8772 7296 8892 7324
rect 8665 7287 8723 7293
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 4580 7228 4905 7256
rect 4580 7216 4586 7228
rect 4893 7225 4905 7228
rect 4939 7225 4951 7259
rect 4893 7219 4951 7225
rect 6454 7216 6460 7268
rect 6512 7256 6518 7268
rect 8864 7265 8892 7296
rect 9858 7284 9864 7336
rect 9916 7284 9922 7336
rect 7377 7259 7435 7265
rect 7377 7256 7389 7259
rect 6512 7228 7389 7256
rect 6512 7216 6518 7228
rect 7377 7225 7389 7228
rect 7423 7225 7435 7259
rect 7377 7219 7435 7225
rect 8849 7259 8907 7265
rect 8849 7225 8861 7259
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 9180 7228 9505 7256
rect 9180 7216 9186 7228
rect 9493 7225 9505 7228
rect 9539 7225 9551 7259
rect 9493 7219 9551 7225
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4304 7160 4721 7188
rect 4304 7148 4310 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 1104 7098 10856 7120
rect 1104 7046 2169 7098
rect 2221 7046 2233 7098
rect 2285 7046 2297 7098
rect 2349 7046 2361 7098
rect 2413 7046 2425 7098
rect 2477 7046 4607 7098
rect 4659 7046 4671 7098
rect 4723 7046 4735 7098
rect 4787 7046 4799 7098
rect 4851 7046 4863 7098
rect 4915 7046 7045 7098
rect 7097 7046 7109 7098
rect 7161 7046 7173 7098
rect 7225 7046 7237 7098
rect 7289 7046 7301 7098
rect 7353 7046 9483 7098
rect 9535 7046 9547 7098
rect 9599 7046 9611 7098
rect 9663 7046 9675 7098
rect 9727 7046 9739 7098
rect 9791 7046 10856 7098
rect 1104 7024 10856 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 5810 6984 5816 6996
rect 2004 6956 5816 6984
rect 2004 6944 2010 6956
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8628 6956 8953 6984
rect 8628 6944 8634 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 6457 6919 6515 6925
rect 6457 6916 6469 6919
rect 6052 6888 6469 6916
rect 6052 6876 6058 6888
rect 6457 6885 6469 6888
rect 6503 6885 6515 6919
rect 9858 6916 9864 6928
rect 6457 6879 6515 6885
rect 8772 6888 9864 6916
rect 1854 6808 1860 6860
rect 1912 6848 1918 6860
rect 2222 6848 2228 6860
rect 1912 6820 2228 6848
rect 1912 6808 1918 6820
rect 2222 6808 2228 6820
rect 2280 6848 2286 6860
rect 6012 6848 6040 6876
rect 2280 6820 5488 6848
rect 2280 6808 2286 6820
rect 1762 6672 1768 6724
rect 1820 6712 1826 6724
rect 5460 6712 5488 6820
rect 5552 6820 6040 6848
rect 6472 6848 6500 6879
rect 6472 6820 6960 6848
rect 5552 6789 5580 6820
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 6043 6752 6101 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6089 6749 6101 6752
rect 6135 6780 6147 6783
rect 6730 6780 6736 6792
rect 6135 6752 6736 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 6932 6789 6960 6820
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 8772 6780 8800 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 8904 6820 9321 6848
rect 8904 6808 8910 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 10042 6808 10048 6860
rect 10100 6848 10106 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10100 6820 10333 6848
rect 10100 6808 10106 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 6963 6752 8800 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 6178 6712 6184 6724
rect 1820 6684 2774 6712
rect 5460 6684 6184 6712
rect 1820 6672 1826 6684
rect 2746 6644 2774 6684
rect 6178 6672 6184 6684
rect 6236 6712 6242 6724
rect 7285 6715 7343 6721
rect 6236 6684 6592 6712
rect 6236 6672 6242 6684
rect 6564 6656 6592 6684
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 7374 6712 7380 6724
rect 7331 6684 7380 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 7374 6672 7380 6684
rect 7432 6712 7438 6724
rect 9416 6712 9444 6743
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 10008 6752 10149 6780
rect 10008 6740 10014 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 7432 6684 9444 6712
rect 7432 6672 7438 6684
rect 5902 6644 5908 6656
rect 2746 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 9272 6616 9689 6644
rect 9272 6604 9278 6616
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 9677 6607 9735 6613
rect 1104 6554 10856 6576
rect 1104 6502 2829 6554
rect 2881 6502 2893 6554
rect 2945 6502 2957 6554
rect 3009 6502 3021 6554
rect 3073 6502 3085 6554
rect 3137 6502 5267 6554
rect 5319 6502 5331 6554
rect 5383 6502 5395 6554
rect 5447 6502 5459 6554
rect 5511 6502 5523 6554
rect 5575 6502 7705 6554
rect 7757 6502 7769 6554
rect 7821 6502 7833 6554
rect 7885 6502 7897 6554
rect 7949 6502 7961 6554
rect 8013 6502 10143 6554
rect 10195 6502 10207 6554
rect 10259 6502 10271 6554
rect 10323 6502 10335 6554
rect 10387 6502 10399 6554
rect 10451 6502 10856 6554
rect 1104 6480 10856 6502
rect 2774 6440 2780 6452
rect 2424 6412 2780 6440
rect 2222 6332 2228 6384
rect 2280 6332 2286 6384
rect 2424 6381 2452 6412
rect 2774 6400 2780 6412
rect 2832 6440 2838 6452
rect 3602 6440 3608 6452
rect 2832 6412 3608 6440
rect 2832 6400 2838 6412
rect 3602 6400 3608 6412
rect 3660 6440 3666 6452
rect 4357 6443 4415 6449
rect 4357 6440 4369 6443
rect 3660 6412 4369 6440
rect 3660 6400 3666 6412
rect 4357 6409 4369 6412
rect 4403 6409 4415 6443
rect 4357 6403 4415 6409
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9122 6440 9128 6452
rect 9079 6412 9128 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 2409 6375 2467 6381
rect 2409 6341 2421 6375
rect 2455 6341 2467 6375
rect 2409 6335 2467 6341
rect 4154 6332 4160 6384
rect 4212 6332 4218 6384
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 9861 6375 9919 6381
rect 9861 6372 9873 6375
rect 6788 6344 9873 6372
rect 6788 6332 6794 6344
rect 9861 6341 9873 6344
rect 9907 6341 9919 6375
rect 9861 6335 9919 6341
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3694 6304 3700 6316
rect 3108 6276 3700 6304
rect 3108 6264 3114 6276
rect 3694 6264 3700 6276
rect 3752 6304 3758 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 3752 6276 5365 6304
rect 3752 6264 3758 6276
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8812 6276 8861 6304
rect 8812 6264 8818 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 10410 6264 10416 6316
rect 10468 6264 10474 6316
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5132 6208 5273 6236
rect 5132 6196 5138 6208
rect 5261 6205 5273 6208
rect 5307 6205 5319 6239
rect 5261 6199 5319 6205
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8444 6208 9137 6236
rect 8444 6196 8450 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 10042 6236 10048 6248
rect 9723 6208 10048 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 3418 6168 3424 6180
rect 1627 6140 3424 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 9585 6171 9643 6177
rect 9585 6168 9597 6171
rect 9456 6140 9597 6168
rect 9456 6128 9462 6140
rect 9585 6137 9597 6140
rect 9631 6137 9643 6171
rect 9585 6131 9643 6137
rect 2038 6060 2044 6112
rect 2096 6060 2102 6112
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 4430 6100 4436 6112
rect 4387 6072 4436 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4522 6060 4528 6112
rect 4580 6060 4586 6112
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 4982 6100 4988 6112
rect 4847 6072 4988 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5442 6060 5448 6112
rect 5500 6060 5506 6112
rect 1104 6010 10856 6032
rect 1104 5958 2169 6010
rect 2221 5958 2233 6010
rect 2285 5958 2297 6010
rect 2349 5958 2361 6010
rect 2413 5958 2425 6010
rect 2477 5958 4607 6010
rect 4659 5958 4671 6010
rect 4723 5958 4735 6010
rect 4787 5958 4799 6010
rect 4851 5958 4863 6010
rect 4915 5958 7045 6010
rect 7097 5958 7109 6010
rect 7161 5958 7173 6010
rect 7225 5958 7237 6010
rect 7289 5958 7301 6010
rect 7353 5958 9483 6010
rect 9535 5958 9547 6010
rect 9599 5958 9611 6010
rect 9663 5958 9675 6010
rect 9727 5958 9739 6010
rect 9791 5958 10856 6010
rect 1104 5936 10856 5958
rect 5166 5896 5172 5908
rect 3528 5868 5172 5896
rect 1946 5788 1952 5840
rect 2004 5828 2010 5840
rect 3142 5828 3148 5840
rect 2004 5800 2360 5828
rect 2004 5788 2010 5800
rect 2038 5720 2044 5772
rect 2096 5720 2102 5772
rect 2332 5701 2360 5800
rect 2792 5800 3148 5828
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2792 5769 2820 5800
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 2685 5763 2743 5769
rect 2685 5760 2697 5763
rect 2648 5732 2697 5760
rect 2648 5720 2654 5732
rect 2685 5729 2697 5732
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 2958 5760 2964 5772
rect 2915 5732 2964 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3234 5760 3240 5772
rect 3099 5732 3240 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3528 5760 3556 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7282 5896 7288 5908
rect 6604 5868 7288 5896
rect 6604 5856 6610 5868
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 8570 5896 8576 5908
rect 7708 5868 8576 5896
rect 7708 5856 7714 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 8996 5868 9413 5896
rect 8996 5856 9002 5868
rect 9401 5865 9413 5868
rect 9447 5865 9459 5899
rect 9401 5859 9459 5865
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 5718 5828 5724 5840
rect 3844 5800 4384 5828
rect 3844 5788 3850 5800
rect 4154 5760 4160 5772
rect 3344 5732 3556 5760
rect 3804 5732 4160 5760
rect 3344 5704 3372 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2317 5695 2375 5701
rect 1627 5664 2268 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1670 5584 1676 5636
rect 1728 5584 1734 5636
rect 1762 5584 1768 5636
rect 1820 5584 1826 5636
rect 1903 5627 1961 5633
rect 1903 5593 1915 5627
rect 1949 5624 1961 5627
rect 1949 5596 2176 5624
rect 1949 5593 1961 5596
rect 1903 5587 1961 5593
rect 1394 5516 1400 5568
rect 1452 5516 1458 5568
rect 2148 5565 2176 5596
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5525 2191 5559
rect 2240 5556 2268 5664
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 3145 5695 3203 5701
rect 2455 5664 2820 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 2332 5624 2360 5655
rect 2792 5636 2820 5664
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3326 5692 3332 5704
rect 3191 5664 3332 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3418 5652 3424 5704
rect 3476 5652 3482 5704
rect 3804 5701 3832 5732
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 4356 5769 4384 5800
rect 4724 5800 5724 5828
rect 4724 5769 4752 5800
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 5902 5788 5908 5840
rect 5960 5828 5966 5840
rect 6914 5828 6920 5840
rect 5960 5800 6920 5828
rect 5960 5788 5966 5800
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 9950 5788 9956 5840
rect 10008 5788 10014 5840
rect 10321 5831 10379 5837
rect 10321 5828 10333 5831
rect 10152 5800 10333 5828
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 4709 5763 4767 5769
rect 4709 5729 4721 5763
rect 4755 5729 4767 5763
rect 4709 5723 4767 5729
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 4982 5760 4988 5772
rect 4847 5732 4988 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5626 5760 5632 5772
rect 5184 5732 5632 5760
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 2682 5624 2688 5636
rect 2332 5596 2688 5624
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 2774 5584 2780 5636
rect 2832 5584 2838 5636
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 3108 5596 3249 5624
rect 3108 5584 3114 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3436 5624 3464 5652
rect 4080 5624 4108 5655
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 5184 5701 5212 5732
rect 5626 5720 5632 5732
rect 5684 5760 5690 5772
rect 6638 5760 6644 5772
rect 5684 5732 6644 5760
rect 5684 5720 5690 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 10152 5769 10180 5800
rect 10321 5797 10333 5800
rect 10367 5797 10379 5831
rect 10321 5791 10379 5797
rect 7929 5763 7987 5769
rect 7929 5760 7941 5763
rect 6748 5732 7941 5760
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4580 5664 4905 5692
rect 4580 5652 4586 5664
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 6748 5701 6776 5732
rect 7929 5729 7941 5732
rect 7975 5729 7987 5763
rect 10137 5763 10195 5769
rect 7929 5723 7987 5729
rect 8864 5732 9996 5760
rect 8864 5704 8892 5732
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 3436 5596 4108 5624
rect 4249 5627 4307 5633
rect 3237 5587 3295 5593
rect 4249 5593 4261 5627
rect 4295 5624 4307 5627
rect 5552 5624 5580 5655
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7190 5652 7196 5704
rect 7248 5652 7254 5704
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8846 5692 8852 5704
rect 8343 5664 8852 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 4295 5596 5580 5624
rect 6825 5627 6883 5633
rect 4295 5593 4307 5596
rect 4249 5587 4307 5593
rect 6825 5593 6837 5627
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 7055 5627 7113 5633
rect 7055 5593 7067 5627
rect 7101 5624 7113 5627
rect 7466 5624 7472 5636
rect 7101 5596 7472 5624
rect 7101 5593 7113 5596
rect 7055 5587 7113 5593
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2240 5528 2881 5556
rect 2133 5519 2191 5525
rect 2869 5525 2881 5528
rect 2915 5525 2927 5559
rect 2869 5519 2927 5525
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 3200 5528 3617 5556
rect 3200 5516 3206 5528
rect 3605 5525 3617 5528
rect 3651 5556 3663 5559
rect 3786 5556 3792 5568
rect 3651 5528 3792 5556
rect 3651 5525 3663 5528
rect 3605 5519 3663 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 4430 5556 4436 5568
rect 3927 5528 4436 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5684 5528 5733 5556
rect 5684 5516 5690 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 5721 5519 5779 5525
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 6512 5528 6561 5556
rect 6512 5516 6518 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 6840 5556 6868 5587
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 7852 5624 7880 5655
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 8938 5652 8944 5704
rect 8996 5652 9002 5704
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 9968 5701 9996 5732
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 9456 5664 9597 5692
rect 9456 5652 9462 5664
rect 9585 5661 9597 5664
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 8018 5624 8024 5636
rect 7852 5596 8024 5624
rect 8018 5584 8024 5596
rect 8076 5624 8082 5636
rect 8113 5627 8171 5633
rect 8113 5624 8125 5627
rect 8076 5596 8125 5624
rect 8076 5584 8082 5596
rect 8113 5593 8125 5596
rect 8159 5624 8171 5627
rect 8389 5627 8447 5633
rect 8389 5624 8401 5627
rect 8159 5596 8401 5624
rect 8159 5593 8171 5596
rect 8113 5587 8171 5593
rect 8389 5593 8401 5596
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 7558 5556 7564 5568
rect 6840 5528 7564 5556
rect 6549 5519 6607 5525
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7745 5559 7803 5565
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 8202 5556 8208 5568
rect 7791 5528 8208 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8404 5556 8432 5587
rect 8570 5584 8576 5636
rect 8628 5584 8634 5636
rect 10152 5624 10180 5723
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 10594 5692 10600 5704
rect 10551 5664 10600 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 8680 5596 10180 5624
rect 8680 5556 8708 5596
rect 8404 5528 8708 5556
rect 8754 5516 8760 5568
rect 8812 5516 8818 5568
rect 1104 5466 10856 5488
rect 1104 5414 2829 5466
rect 2881 5414 2893 5466
rect 2945 5414 2957 5466
rect 3009 5414 3021 5466
rect 3073 5414 3085 5466
rect 3137 5414 5267 5466
rect 5319 5414 5331 5466
rect 5383 5414 5395 5466
rect 5447 5414 5459 5466
rect 5511 5414 5523 5466
rect 5575 5414 7705 5466
rect 7757 5414 7769 5466
rect 7821 5414 7833 5466
rect 7885 5414 7897 5466
rect 7949 5414 7961 5466
rect 8013 5414 10143 5466
rect 10195 5414 10207 5466
rect 10259 5414 10271 5466
rect 10323 5414 10335 5466
rect 10387 5414 10399 5466
rect 10451 5414 10856 5466
rect 1104 5392 10856 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1489 5355 1547 5361
rect 1489 5352 1501 5355
rect 1360 5324 1501 5352
rect 1360 5312 1366 5324
rect 1489 5321 1501 5324
rect 1535 5321 1547 5355
rect 1489 5315 1547 5321
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 2317 5355 2375 5361
rect 2317 5352 2329 5355
rect 1728 5324 2329 5352
rect 1728 5312 1734 5324
rect 2317 5321 2329 5324
rect 2363 5321 2375 5355
rect 2317 5315 2375 5321
rect 3602 5312 3608 5364
rect 3660 5312 3666 5364
rect 4449 5355 4507 5361
rect 4449 5352 4461 5355
rect 3804 5324 4461 5352
rect 1394 5244 1400 5296
rect 1452 5284 1458 5296
rect 3804 5293 3832 5324
rect 4449 5321 4461 5324
rect 4495 5321 4507 5355
rect 4449 5315 4507 5321
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 5166 5352 5172 5364
rect 4663 5324 5172 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 7190 5352 7196 5364
rect 6779 5324 7196 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 7466 5312 7472 5364
rect 7524 5312 7530 5364
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 1452 5256 1992 5284
rect 1452 5244 1458 5256
rect 1964 5225 1992 5256
rect 3528 5256 3801 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1949 5219 2007 5225
rect 1719 5188 1808 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1780 5089 1808 5188
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 3234 5216 3240 5228
rect 2731 5188 3240 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 3528 5225 3556 5256
rect 3789 5253 3801 5256
rect 3835 5253 3847 5287
rect 3789 5247 3847 5253
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4249 5287 4307 5293
rect 4249 5284 4261 5287
rect 4212 5256 4261 5284
rect 4212 5244 4218 5256
rect 4249 5253 4261 5256
rect 4295 5253 4307 5287
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 4249 5247 4307 5253
rect 7024 5256 7849 5284
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3476 5188 3525 5216
rect 3476 5176 3482 5188
rect 3513 5185 3525 5188
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4172 5216 4200 5244
rect 4111 5188 4200 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 2498 5108 2504 5160
rect 2556 5148 2562 5160
rect 2593 5151 2651 5157
rect 2593 5148 2605 5151
rect 2556 5120 2605 5148
rect 2556 5108 2562 5120
rect 2593 5117 2605 5120
rect 2639 5148 2651 5151
rect 3712 5148 3740 5176
rect 2639 5120 3740 5148
rect 3988 5148 4016 5179
rect 6454 5176 6460 5228
rect 6512 5176 6518 5228
rect 7024 5225 7052 5256
rect 7837 5253 7849 5256
rect 7883 5284 7895 5287
rect 8202 5284 8208 5296
rect 7883 5256 8208 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 7466 5216 7472 5228
rect 7331 5188 7472 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7650 5176 7656 5228
rect 7708 5176 7714 5228
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8386 5216 8392 5228
rect 8343 5188 8392 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8628 5188 9045 5216
rect 8628 5176 8634 5188
rect 9033 5185 9045 5188
rect 9079 5216 9091 5219
rect 9306 5216 9312 5228
rect 9079 5188 9312 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9306 5176 9312 5188
rect 9364 5216 9370 5228
rect 10336 5216 10364 5315
rect 9364 5188 10364 5216
rect 9364 5176 9370 5188
rect 10502 5176 10508 5228
rect 10560 5176 10566 5228
rect 4430 5148 4436 5160
rect 3988 5120 4436 5148
rect 2639 5117 2651 5120
rect 2593 5111 2651 5117
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6788 5120 6929 5148
rect 6788 5108 6794 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5049 1823 5083
rect 1765 5043 1823 5049
rect 3234 5040 3240 5092
rect 3292 5080 3298 5092
rect 3789 5083 3847 5089
rect 3789 5080 3801 5083
rect 3292 5052 3801 5080
rect 3292 5040 3298 5052
rect 3789 5049 3801 5052
rect 3835 5049 3847 5083
rect 3789 5043 3847 5049
rect 2685 5015 2743 5021
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 3326 5012 3332 5024
rect 2731 4984 3332 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 4448 5021 4476 5108
rect 6641 5083 6699 5089
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 7392 5080 7420 5111
rect 8754 5080 8760 5092
rect 6687 5052 6960 5080
rect 7392 5052 8760 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 6932 5024 6960 5052
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 9306 5080 9312 5092
rect 8904 5052 9312 5080
rect 8904 5040 8910 5052
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 4981 4491 5015
rect 4433 4975 4491 4981
rect 6914 4972 6920 5024
rect 6972 4972 6978 5024
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 7650 5012 7656 5024
rect 7340 4984 7656 5012
rect 7340 4972 7346 4984
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 1104 4922 10856 4944
rect 1104 4870 2169 4922
rect 2221 4870 2233 4922
rect 2285 4870 2297 4922
rect 2349 4870 2361 4922
rect 2413 4870 2425 4922
rect 2477 4870 4607 4922
rect 4659 4870 4671 4922
rect 4723 4870 4735 4922
rect 4787 4870 4799 4922
rect 4851 4870 4863 4922
rect 4915 4870 7045 4922
rect 7097 4870 7109 4922
rect 7161 4870 7173 4922
rect 7225 4870 7237 4922
rect 7289 4870 7301 4922
rect 7353 4870 9483 4922
rect 9535 4870 9547 4922
rect 9599 4870 9611 4922
rect 9663 4870 9675 4922
rect 9727 4870 9739 4922
rect 9791 4870 10856 4922
rect 1104 4848 10856 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 2498 4808 2504 4820
rect 1627 4780 2504 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5868 4780 6009 4808
rect 5868 4768 5874 4780
rect 5997 4777 6009 4780
rect 6043 4808 6055 4811
rect 6730 4808 6736 4820
rect 6043 4780 6736 4808
rect 6043 4777 6055 4780
rect 5997 4771 6055 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 8021 4811 8079 4817
rect 8021 4808 8033 4811
rect 7616 4780 8033 4808
rect 7616 4768 7622 4780
rect 8021 4777 8033 4780
rect 8067 4777 8079 4811
rect 8021 4771 8079 4777
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8128 4712 9045 4740
rect 6638 4632 6644 4684
rect 6696 4632 6702 4684
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 7374 4672 7380 4684
rect 7331 4644 7380 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6454 4604 6460 4616
rect 6135 4576 6460 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 6917 4607 6975 4613
rect 6917 4604 6929 4607
rect 6880 4576 6929 4604
rect 6880 4564 6886 4576
rect 6917 4573 6929 4576
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4604 7987 4607
rect 8018 4604 8024 4616
rect 7975 4576 8024 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8128 4613 8156 4712
rect 9033 4709 9045 4712
rect 9079 4709 9091 4743
rect 9033 4703 9091 4709
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8294 4672 8300 4684
rect 8251 4644 8300 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 8938 4672 8944 4684
rect 8803 4644 8944 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 9493 4675 9551 4681
rect 9493 4672 9505 4675
rect 9364 4644 9505 4672
rect 9364 4632 9370 4644
rect 9493 4641 9505 4644
rect 9539 4641 9551 4675
rect 9493 4635 9551 4641
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9030 4604 9036 4616
rect 8711 4576 9036 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8294 4536 8300 4548
rect 7760 4508 8300 4536
rect 7760 4477 7788 4508
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4437 7803 4471
rect 7745 4431 7803 4437
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 8404 4468 8432 4567
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 8260 4440 8432 4468
rect 8260 4428 8266 4440
rect 1104 4378 10856 4400
rect 1104 4326 2829 4378
rect 2881 4326 2893 4378
rect 2945 4326 2957 4378
rect 3009 4326 3021 4378
rect 3073 4326 3085 4378
rect 3137 4326 5267 4378
rect 5319 4326 5331 4378
rect 5383 4326 5395 4378
rect 5447 4326 5459 4378
rect 5511 4326 5523 4378
rect 5575 4326 7705 4378
rect 7757 4326 7769 4378
rect 7821 4326 7833 4378
rect 7885 4326 7897 4378
rect 7949 4326 7961 4378
rect 8013 4326 10143 4378
rect 10195 4326 10207 4378
rect 10259 4326 10271 4378
rect 10323 4326 10335 4378
rect 10387 4326 10399 4378
rect 10451 4326 10856 4378
rect 1104 4304 10856 4326
rect 5505 4199 5563 4205
rect 5505 4196 5517 4199
rect 4264 4168 5517 4196
rect 4264 4137 4292 4168
rect 5505 4165 5517 4168
rect 5551 4196 5563 4199
rect 5551 4168 5672 4196
rect 5551 4165 5563 4168
rect 5505 4159 5563 4165
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4264 4060 4292 4091
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4396 4100 4445 4128
rect 4396 4088 4402 4100
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 5644 4128 5672 4168
rect 5718 4156 5724 4208
rect 5776 4196 5782 4208
rect 5776 4168 6132 4196
rect 5776 4156 5782 4168
rect 6104 4137 6132 4168
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 6788 4168 7328 4196
rect 6788 4156 6794 4168
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5644 4100 5825 4128
rect 4433 4091 4491 4097
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4097 6147 4131
rect 7300 4128 7328 4168
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 7432 4168 7880 4196
rect 7432 4156 7438 4168
rect 7852 4137 7880 4168
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7300 4100 7665 4128
rect 6089 4091 6147 4097
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 4264 4032 4476 4060
rect 4448 4004 4476 4032
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5261 4063 5319 4069
rect 5261 4060 5273 4063
rect 5132 4032 5273 4060
rect 5132 4020 5138 4032
rect 5261 4029 5273 4032
rect 5307 4029 5319 4063
rect 5261 4023 5319 4029
rect 4430 3952 4436 4004
rect 4488 3952 4494 4004
rect 5276 3992 5304 4023
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 6012 4060 6040 4091
rect 8938 4088 8944 4140
rect 8996 4088 9002 4140
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 9858 4128 9864 4140
rect 9815 4100 9864 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 5684 4032 6040 4060
rect 7561 4063 7619 4069
rect 5684 4020 5690 4032
rect 7561 4029 7573 4063
rect 7607 4060 7619 4063
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 7607 4032 8217 4060
rect 7607 4029 7619 4032
rect 7561 4023 7619 4029
rect 8205 4029 8217 4032
rect 8251 4060 8263 4063
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8251 4032 8677 4060
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 8665 4029 8677 4032
rect 8711 4060 8723 4063
rect 8846 4060 8852 4072
rect 8711 4032 8852 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 5276 3964 7113 3992
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 7101 3955 7159 3961
rect 4338 3884 4344 3936
rect 4396 3884 4402 3936
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 4801 3927 4859 3933
rect 4801 3924 4813 3927
rect 4580 3896 4813 3924
rect 4580 3884 4586 3896
rect 4801 3893 4813 3896
rect 4847 3893 4859 3927
rect 4801 3887 4859 3893
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 5040 3896 5365 3924
rect 5040 3884 5046 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5353 3887 5411 3893
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3924 5595 3927
rect 5626 3924 5632 3936
rect 5583 3896 5632 3924
rect 5583 3893 5595 3896
rect 5537 3887 5595 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9456 3896 9597 3924
rect 9456 3884 9462 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9585 3887 9643 3893
rect 1104 3834 10856 3856
rect 1104 3782 2169 3834
rect 2221 3782 2233 3834
rect 2285 3782 2297 3834
rect 2349 3782 2361 3834
rect 2413 3782 2425 3834
rect 2477 3782 4607 3834
rect 4659 3782 4671 3834
rect 4723 3782 4735 3834
rect 4787 3782 4799 3834
rect 4851 3782 4863 3834
rect 4915 3782 7045 3834
rect 7097 3782 7109 3834
rect 7161 3782 7173 3834
rect 7225 3782 7237 3834
rect 7289 3782 7301 3834
rect 7353 3782 9483 3834
rect 9535 3782 9547 3834
rect 9599 3782 9611 3834
rect 9663 3782 9675 3834
rect 9727 3782 9739 3834
rect 9791 3782 10856 3834
rect 1104 3760 10856 3782
rect 2682 3680 2688 3732
rect 2740 3720 2746 3732
rect 4614 3720 4620 3732
rect 2740 3692 4620 3720
rect 2740 3680 2746 3692
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 2832 3624 3188 3652
rect 2832 3612 2838 3624
rect 842 3544 848 3596
rect 900 3584 906 3596
rect 1489 3587 1547 3593
rect 1489 3584 1501 3587
rect 900 3556 1501 3584
rect 900 3544 906 3556
rect 1489 3553 1501 3556
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 3160 3593 3188 3624
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 4724 3652 4752 3683
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 9122 3720 9128 3732
rect 6696 3692 9128 3720
rect 6696 3680 6702 3692
rect 9122 3680 9128 3692
rect 9180 3720 9186 3732
rect 10042 3720 10048 3732
rect 9180 3692 10048 3720
rect 9180 3680 9186 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 4580 3624 4752 3652
rect 7469 3655 7527 3661
rect 4580 3612 4586 3624
rect 7469 3621 7481 3655
rect 7515 3652 7527 3655
rect 7561 3655 7619 3661
rect 7561 3652 7573 3655
rect 7515 3624 7573 3652
rect 7515 3621 7527 3624
rect 7469 3615 7527 3621
rect 7561 3621 7573 3624
rect 7607 3621 7619 3655
rect 7561 3615 7619 3621
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 8444 3624 10272 3652
rect 8444 3612 8450 3624
rect 2501 3587 2559 3593
rect 1820 3556 2176 3584
rect 1820 3544 1826 3556
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 2148 3516 2176 3556
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 3145 3587 3203 3593
rect 2547 3556 3096 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2148 3488 2605 3516
rect 2593 3485 2605 3488
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2682 3476 2688 3528
rect 2740 3476 2746 3528
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 3068 3448 3096 3556
rect 3145 3553 3157 3587
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 3510 3544 3516 3596
rect 3568 3544 3574 3596
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4212 3556 4384 3584
rect 4212 3544 4218 3556
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3326 3516 3332 3528
rect 3283 3488 3332 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 4356 3525 4384 3556
rect 4614 3544 4620 3596
rect 4672 3584 4678 3596
rect 5166 3584 5172 3596
rect 4672 3556 5172 3584
rect 4672 3544 4678 3556
rect 5166 3544 5172 3556
rect 5224 3584 5230 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5224 3556 5457 3584
rect 5224 3544 5230 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5583 3556 5917 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7374 3584 7380 3596
rect 6963 3556 7380 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 7852 3556 8769 3584
rect 4341 3519 4399 3525
rect 3988 3488 4292 3516
rect 3418 3448 3424 3460
rect 3068 3420 3424 3448
rect 3418 3408 3424 3420
rect 3476 3408 3482 3460
rect 3988 3457 4016 3488
rect 3605 3451 3663 3457
rect 3605 3417 3617 3451
rect 3651 3448 3663 3451
rect 3973 3451 4031 3457
rect 3973 3448 3985 3451
rect 3651 3420 3985 3448
rect 3651 3417 3663 3420
rect 3605 3411 3663 3417
rect 3973 3417 3985 3420
rect 4019 3417 4031 3451
rect 3973 3411 4031 3417
rect 4157 3451 4215 3457
rect 4157 3417 4169 3451
rect 4203 3417 4215 3451
rect 4264 3448 4292 3488
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4448 3448 4476 3479
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4580 3488 4721 3516
rect 4580 3476 4586 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5718 3516 5724 3528
rect 5132 3488 5724 3516
rect 5132 3476 5138 3488
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 4264 3420 4476 3448
rect 5000 3448 5028 3476
rect 5828 3448 5856 3479
rect 5000 3420 5856 3448
rect 6012 3448 6040 3479
rect 7558 3476 7564 3528
rect 7616 3476 7622 3528
rect 7852 3525 7880 3556
rect 8757 3553 8769 3556
rect 8803 3553 8815 3587
rect 8757 3547 8815 3553
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 10244 3593 10272 3624
rect 10229 3587 10287 3593
rect 8904 3556 9812 3584
rect 8904 3544 8910 3556
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8067 3488 8248 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 6638 3448 6644 3460
rect 6012 3420 6644 3448
rect 4157 3411 4215 3417
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 2280 3352 2329 3380
rect 2280 3340 2286 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 3234 3380 3240 3392
rect 3007 3352 3240 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 3234 3340 3240 3352
rect 3292 3340 3298 3392
rect 4172 3380 4200 3411
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 7576 3448 7604 3476
rect 7116 3420 7604 3448
rect 7116 3392 7144 3420
rect 4430 3380 4436 3392
rect 4172 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 5031 3352 5089 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5077 3349 5089 3352
rect 5123 3349 5135 3383
rect 5077 3343 5135 3349
rect 5718 3340 5724 3392
rect 5776 3340 5782 3392
rect 7006 3340 7012 3392
rect 7064 3340 7070 3392
rect 7098 3340 7104 3392
rect 7156 3340 7162 3392
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7616 3352 7757 3380
rect 7616 3340 7622 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 8220 3380 8248 3488
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8478 3476 8484 3528
rect 8536 3476 8542 3528
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 8588 3448 8616 3479
rect 8938 3476 8944 3528
rect 8996 3476 9002 3528
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 9306 3476 9312 3528
rect 9364 3476 9370 3528
rect 9674 3476 9680 3528
rect 9732 3476 9738 3528
rect 9784 3516 9812 3556
rect 10229 3553 10241 3587
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 9870 3519 9928 3525
rect 9870 3516 9882 3519
rect 9784 3488 9882 3516
rect 9870 3485 9882 3488
rect 9916 3485 9928 3519
rect 9870 3479 9928 3485
rect 9398 3448 9404 3460
rect 8588 3420 9404 3448
rect 9398 3408 9404 3420
rect 9456 3408 9462 3460
rect 8938 3380 8944 3392
rect 8220 3352 8944 3380
rect 7745 3343 7803 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 1104 3290 10856 3312
rect 1104 3238 2829 3290
rect 2881 3238 2893 3290
rect 2945 3238 2957 3290
rect 3009 3238 3021 3290
rect 3073 3238 3085 3290
rect 3137 3238 5267 3290
rect 5319 3238 5331 3290
rect 5383 3238 5395 3290
rect 5447 3238 5459 3290
rect 5511 3238 5523 3290
rect 5575 3238 7705 3290
rect 7757 3238 7769 3290
rect 7821 3238 7833 3290
rect 7885 3238 7897 3290
rect 7949 3238 7961 3290
rect 8013 3238 10143 3290
rect 10195 3238 10207 3290
rect 10259 3238 10271 3290
rect 10323 3238 10335 3290
rect 10387 3238 10399 3290
rect 10451 3238 10856 3290
rect 1104 3216 10856 3238
rect 2038 3136 2044 3188
rect 2096 3136 2102 3188
rect 2774 3136 2780 3188
rect 2832 3136 2838 3188
rect 3418 3136 3424 3188
rect 3476 3176 3482 3188
rect 3973 3179 4031 3185
rect 3973 3176 3985 3179
rect 3476 3148 3985 3176
rect 3476 3136 3482 3148
rect 3973 3145 3985 3148
rect 4019 3145 4031 3179
rect 3973 3139 4031 3145
rect 4522 3136 4528 3188
rect 4580 3136 4586 3188
rect 5074 3176 5080 3188
rect 4908 3148 5080 3176
rect 3234 3068 3240 3120
rect 3292 3068 3298 3120
rect 4338 3068 4344 3120
rect 4396 3108 4402 3120
rect 4908 3117 4936 3148
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 5224 3148 5457 3176
rect 5224 3136 5230 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7432 3148 7849 3176
rect 7432 3136 7438 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 8938 3176 8944 3188
rect 8803 3148 8944 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9125 3179 9183 3185
rect 9125 3145 9137 3179
rect 9171 3176 9183 3179
rect 9306 3176 9312 3188
rect 9171 3148 9312 3176
rect 9171 3145 9183 3148
rect 9125 3139 9183 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9582 3176 9588 3188
rect 9416 3148 9588 3176
rect 4677 3111 4735 3117
rect 4677 3108 4689 3111
rect 4396 3080 4689 3108
rect 4396 3068 4402 3080
rect 4677 3077 4689 3080
rect 4723 3077 4735 3111
rect 4677 3071 4735 3077
rect 4893 3111 4951 3117
rect 4893 3077 4905 3111
rect 4939 3077 4951 3111
rect 5810 3108 5816 3120
rect 4893 3071 4951 3077
rect 5092 3080 5816 3108
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3252 3040 3280 3068
rect 4062 3040 4068 3052
rect 3007 3012 3280 3040
rect 3896 3012 4068 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3896 2972 3924 3012
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4982 3040 4988 3052
rect 4295 3012 4988 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5092 3049 5120 3080
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 3283 2944 3924 2972
rect 3973 2975 4031 2981
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4154 2972 4160 2984
rect 4019 2944 4160 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4154 2932 4160 2944
rect 4212 2972 4218 2984
rect 5276 2972 5304 3003
rect 4212 2944 5304 2972
rect 4212 2932 4218 2944
rect 3145 2907 3203 2913
rect 3145 2873 3157 2907
rect 3191 2904 3203 2907
rect 3326 2904 3332 2916
rect 3191 2876 3332 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 3326 2864 3332 2876
rect 3384 2904 3390 2916
rect 4338 2904 4344 2916
rect 3384 2876 4344 2904
rect 3384 2864 3390 2876
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 5368 2904 5396 3080
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 7466 3108 7472 3120
rect 7208 3080 7472 3108
rect 7208 3049 7236 3080
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 8662 3108 8668 3120
rect 7852 3080 8668 3108
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 7852 3049 7880 3080
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9416 3108 9444 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9732 3148 9873 3176
rect 9732 3136 9738 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 8864 3080 9444 3108
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2972 7527 2975
rect 7852 2972 7880 3003
rect 7515 2944 7880 2972
rect 8036 2972 8064 3003
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8536 3012 8769 3040
rect 8536 3000 8542 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8386 2972 8392 2984
rect 8036 2944 8392 2972
rect 7515 2941 7527 2944
rect 7469 2935 7527 2941
rect 4632 2876 5396 2904
rect 7377 2907 7435 2913
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4632 2836 4660 2876
rect 7377 2873 7389 2907
rect 7423 2904 7435 2907
rect 8036 2904 8064 2944
rect 8386 2932 8392 2944
rect 8444 2972 8450 2984
rect 8864 2972 8892 3080
rect 9490 3068 9496 3120
rect 9548 3108 9554 3120
rect 9950 3108 9956 3120
rect 9548 3080 9956 3108
rect 9548 3068 9554 3080
rect 9950 3068 9956 3080
rect 10008 3108 10014 3120
rect 10008 3080 10456 3108
rect 10008 3068 10014 3080
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9398 3040 9404 3052
rect 8987 3012 9404 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9398 3000 9404 3012
rect 9456 3040 9462 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9456 3012 9689 3040
rect 9456 3000 9462 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 9858 3000 9864 3052
rect 9916 3040 9922 3052
rect 10428 3049 10456 3080
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 9916 3012 10241 3040
rect 9916 3000 9922 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 8444 2944 8892 2972
rect 8444 2932 8450 2944
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9548 2944 9597 2972
rect 9548 2932 9554 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 7423 2876 8064 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 9214 2864 9220 2916
rect 9272 2904 9278 2916
rect 9309 2907 9367 2913
rect 9309 2904 9321 2907
rect 9272 2876 9321 2904
rect 9272 2864 9278 2876
rect 9309 2873 9321 2876
rect 9355 2904 9367 2907
rect 9876 2904 9904 3000
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 10183 2944 10333 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 9355 2876 9904 2904
rect 9355 2873 9367 2876
rect 9309 2867 9367 2873
rect 4203 2808 4660 2836
rect 4709 2839 4767 2845
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 5626 2836 5632 2848
rect 4755 2808 5632 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 7745 2839 7803 2845
rect 7745 2805 7757 2839
rect 7791 2836 7803 2839
rect 7834 2836 7840 2848
rect 7791 2808 7840 2836
rect 7791 2805 7803 2808
rect 7745 2799 7803 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 10152 2836 10180 2935
rect 8536 2808 10180 2836
rect 8536 2796 8542 2808
rect 1104 2746 10856 2768
rect 1104 2694 2169 2746
rect 2221 2694 2233 2746
rect 2285 2694 2297 2746
rect 2349 2694 2361 2746
rect 2413 2694 2425 2746
rect 2477 2694 4607 2746
rect 4659 2694 4671 2746
rect 4723 2694 4735 2746
rect 4787 2694 4799 2746
rect 4851 2694 4863 2746
rect 4915 2694 7045 2746
rect 7097 2694 7109 2746
rect 7161 2694 7173 2746
rect 7225 2694 7237 2746
rect 7289 2694 7301 2746
rect 7353 2694 9483 2746
rect 9535 2694 9547 2746
rect 9599 2694 9611 2746
rect 9663 2694 9675 2746
rect 9727 2694 9739 2746
rect 9791 2694 10856 2746
rect 1104 2672 10856 2694
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 4430 2592 4436 2644
rect 4488 2632 4494 2644
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4488 2604 4721 2632
rect 4488 2592 4494 2604
rect 4709 2601 4721 2604
rect 4755 2601 4767 2635
rect 4709 2595 4767 2601
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6512 2604 6745 2632
rect 6512 2592 6518 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 9214 2632 9220 2644
rect 8720 2604 9220 2632
rect 8720 2592 8726 2604
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9306 2592 9312 2644
rect 9364 2592 9370 2644
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 9953 2635 10011 2641
rect 9953 2632 9965 2635
rect 9916 2604 9965 2632
rect 9916 2592 9922 2604
rect 9953 2601 9965 2604
rect 9999 2601 10011 2635
rect 9953 2595 10011 2601
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5718 2428 5724 2440
rect 5491 2400 5724 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6972 2400 7205 2428
rect 6972 2388 6978 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8444 2400 8493 2428
rect 8444 2388 8450 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5166 2360 5172 2372
rect 5123 2332 5172 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5166 2320 5172 2332
rect 5224 2320 5230 2372
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 7558 2252 7564 2304
rect 7616 2292 7622 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7616 2264 8033 2292
rect 7616 2252 7622 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 1104 2202 10856 2224
rect 1104 2150 2829 2202
rect 2881 2150 2893 2202
rect 2945 2150 2957 2202
rect 3009 2150 3021 2202
rect 3073 2150 3085 2202
rect 3137 2150 5267 2202
rect 5319 2150 5331 2202
rect 5383 2150 5395 2202
rect 5447 2150 5459 2202
rect 5511 2150 5523 2202
rect 5575 2150 7705 2202
rect 7757 2150 7769 2202
rect 7821 2150 7833 2202
rect 7885 2150 7897 2202
rect 7949 2150 7961 2202
rect 8013 2150 10143 2202
rect 10195 2150 10207 2202
rect 10259 2150 10271 2202
rect 10323 2150 10335 2202
rect 10387 2150 10399 2202
rect 10451 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 7104 11840 7156 11892
rect 8208 11840 8260 11892
rect 2169 11398 2221 11450
rect 2233 11398 2285 11450
rect 2297 11398 2349 11450
rect 2361 11398 2413 11450
rect 2425 11398 2477 11450
rect 4607 11398 4659 11450
rect 4671 11398 4723 11450
rect 4735 11398 4787 11450
rect 4799 11398 4851 11450
rect 4863 11398 4915 11450
rect 7045 11398 7097 11450
rect 7109 11398 7161 11450
rect 7173 11398 7225 11450
rect 7237 11398 7289 11450
rect 7301 11398 7353 11450
rect 9483 11398 9535 11450
rect 9547 11398 9599 11450
rect 9611 11398 9663 11450
rect 9675 11398 9727 11450
rect 9739 11398 9791 11450
rect 5816 11296 5868 11348
rect 4528 11160 4580 11212
rect 3884 11092 3936 11144
rect 5172 11092 5224 11144
rect 7104 11203 7156 11212
rect 7104 11169 7113 11203
rect 7113 11169 7147 11203
rect 7147 11169 7156 11203
rect 7104 11160 7156 11169
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 7472 11092 7524 11144
rect 8208 11092 8260 11144
rect 6460 11067 6512 11076
rect 6460 11033 6469 11067
rect 6469 11033 6503 11067
rect 6503 11033 6512 11067
rect 6460 11024 6512 11033
rect 3884 10956 3936 11008
rect 4252 10956 4304 11008
rect 5080 10956 5132 11008
rect 8300 10956 8352 11008
rect 2829 10854 2881 10906
rect 2893 10854 2945 10906
rect 2957 10854 3009 10906
rect 3021 10854 3073 10906
rect 3085 10854 3137 10906
rect 5267 10854 5319 10906
rect 5331 10854 5383 10906
rect 5395 10854 5447 10906
rect 5459 10854 5511 10906
rect 5523 10854 5575 10906
rect 7705 10854 7757 10906
rect 7769 10854 7821 10906
rect 7833 10854 7885 10906
rect 7897 10854 7949 10906
rect 7961 10854 8013 10906
rect 10143 10854 10195 10906
rect 10207 10854 10259 10906
rect 10271 10854 10323 10906
rect 10335 10854 10387 10906
rect 10399 10854 10451 10906
rect 5080 10795 5132 10804
rect 3424 10684 3476 10736
rect 5080 10761 5107 10795
rect 5107 10761 5132 10795
rect 5080 10752 5132 10761
rect 6460 10752 6512 10804
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2780 10659 2832 10668
rect 2780 10625 2789 10659
rect 2789 10625 2823 10659
rect 2823 10625 2832 10659
rect 2780 10616 2832 10625
rect 3884 10548 3936 10600
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 5264 10727 5316 10736
rect 5264 10693 5273 10727
rect 5273 10693 5307 10727
rect 5307 10693 5316 10727
rect 5264 10684 5316 10693
rect 7104 10752 7156 10804
rect 7472 10752 7524 10804
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 7380 10684 7432 10736
rect 4068 10480 4120 10532
rect 848 10412 900 10464
rect 1676 10412 1728 10464
rect 3240 10412 3292 10464
rect 4436 10412 4488 10464
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7656 10616 7708 10668
rect 8208 10684 8260 10736
rect 8116 10616 8168 10668
rect 7380 10548 7432 10600
rect 8576 10548 8628 10600
rect 8300 10480 8352 10532
rect 5356 10412 5408 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6184 10412 6236 10464
rect 6644 10412 6696 10464
rect 2169 10310 2221 10362
rect 2233 10310 2285 10362
rect 2297 10310 2349 10362
rect 2361 10310 2413 10362
rect 2425 10310 2477 10362
rect 4607 10310 4659 10362
rect 4671 10310 4723 10362
rect 4735 10310 4787 10362
rect 4799 10310 4851 10362
rect 4863 10310 4915 10362
rect 7045 10310 7097 10362
rect 7109 10310 7161 10362
rect 7173 10310 7225 10362
rect 7237 10310 7289 10362
rect 7301 10310 7353 10362
rect 9483 10310 9535 10362
rect 9547 10310 9599 10362
rect 9611 10310 9663 10362
rect 9675 10310 9727 10362
rect 9739 10310 9791 10362
rect 2044 10208 2096 10260
rect 3792 10208 3844 10260
rect 5540 10208 5592 10260
rect 6276 10208 6328 10260
rect 2780 10140 2832 10192
rect 4068 10140 4120 10192
rect 1400 10072 1452 10124
rect 4160 10072 4212 10124
rect 5264 10183 5316 10192
rect 5264 10149 5273 10183
rect 5273 10149 5307 10183
rect 5307 10149 5316 10183
rect 5264 10140 5316 10149
rect 5356 10140 5408 10192
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 3884 10047 3936 10056
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 1768 9979 1820 9988
rect 1768 9945 1777 9979
rect 1777 9945 1811 9979
rect 1811 9945 1820 9979
rect 1768 9936 1820 9945
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 3332 9936 3384 9988
rect 5816 10072 5868 10124
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 7656 10072 7708 10124
rect 7472 10004 7524 10056
rect 4252 9868 4304 9920
rect 4804 9911 4856 9920
rect 4804 9877 4813 9911
rect 4813 9877 4847 9911
rect 4847 9877 4856 9911
rect 4804 9868 4856 9877
rect 5908 9936 5960 9988
rect 6460 9979 6512 9988
rect 6460 9945 6495 9979
rect 6495 9945 6512 9979
rect 6460 9936 6512 9945
rect 8208 10004 8260 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 6828 9868 6880 9920
rect 7012 9868 7064 9920
rect 8300 9868 8352 9920
rect 2829 9766 2881 9818
rect 2893 9766 2945 9818
rect 2957 9766 3009 9818
rect 3021 9766 3073 9818
rect 3085 9766 3137 9818
rect 5267 9766 5319 9818
rect 5331 9766 5383 9818
rect 5395 9766 5447 9818
rect 5459 9766 5511 9818
rect 5523 9766 5575 9818
rect 7705 9766 7757 9818
rect 7769 9766 7821 9818
rect 7833 9766 7885 9818
rect 7897 9766 7949 9818
rect 7961 9766 8013 9818
rect 10143 9766 10195 9818
rect 10207 9766 10259 9818
rect 10271 9766 10323 9818
rect 10335 9766 10387 9818
rect 10399 9766 10451 9818
rect 2136 9664 2188 9716
rect 4620 9664 4672 9716
rect 5632 9664 5684 9716
rect 6276 9664 6328 9716
rect 6460 9664 6512 9716
rect 2504 9596 2556 9648
rect 3792 9639 3844 9648
rect 3792 9605 3801 9639
rect 3801 9605 3835 9639
rect 3835 9605 3844 9639
rect 3792 9596 3844 9605
rect 4804 9596 4856 9648
rect 7012 9639 7064 9648
rect 7012 9605 7021 9639
rect 7021 9605 7055 9639
rect 7055 9605 7064 9639
rect 7012 9596 7064 9605
rect 1952 9528 2004 9580
rect 3240 9528 3292 9580
rect 3424 9528 3476 9580
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 4160 9528 4212 9580
rect 7380 9528 7432 9580
rect 1768 9392 1820 9444
rect 5080 9460 5132 9512
rect 6460 9460 6512 9512
rect 6828 9460 6880 9512
rect 4988 9392 5040 9444
rect 8208 9528 8260 9580
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8576 9460 8628 9512
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 3332 9324 3384 9376
rect 6828 9324 6880 9376
rect 6920 9324 6972 9376
rect 2169 9222 2221 9274
rect 2233 9222 2285 9274
rect 2297 9222 2349 9274
rect 2361 9222 2413 9274
rect 2425 9222 2477 9274
rect 4607 9222 4659 9274
rect 4671 9222 4723 9274
rect 4735 9222 4787 9274
rect 4799 9222 4851 9274
rect 4863 9222 4915 9274
rect 7045 9222 7097 9274
rect 7109 9222 7161 9274
rect 7173 9222 7225 9274
rect 7237 9222 7289 9274
rect 7301 9222 7353 9274
rect 9483 9222 9535 9274
rect 9547 9222 9599 9274
rect 9611 9222 9663 9274
rect 9675 9222 9727 9274
rect 9739 9222 9791 9274
rect 8576 9120 8628 9172
rect 5632 8984 5684 9036
rect 848 8916 900 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9404 8848 9456 8900
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 3240 8780 3292 8832
rect 9036 8780 9088 8832
rect 9864 8780 9916 8832
rect 9956 8780 10008 8832
rect 2829 8678 2881 8730
rect 2893 8678 2945 8730
rect 2957 8678 3009 8730
rect 3021 8678 3073 8730
rect 3085 8678 3137 8730
rect 5267 8678 5319 8730
rect 5331 8678 5383 8730
rect 5395 8678 5447 8730
rect 5459 8678 5511 8730
rect 5523 8678 5575 8730
rect 7705 8678 7757 8730
rect 7769 8678 7821 8730
rect 7833 8678 7885 8730
rect 7897 8678 7949 8730
rect 7961 8678 8013 8730
rect 10143 8678 10195 8730
rect 10207 8678 10259 8730
rect 10271 8678 10323 8730
rect 10335 8678 10387 8730
rect 10399 8678 10451 8730
rect 9128 8576 9180 8628
rect 9956 8551 10008 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1952 8440 2004 8492
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 2596 8440 2648 8492
rect 5172 8440 5224 8492
rect 8668 8440 8720 8492
rect 9956 8517 9965 8551
rect 9965 8517 9999 8551
rect 9999 8517 10008 8551
rect 9956 8508 10008 8517
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9588 8440 9640 8492
rect 9864 8440 9916 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1584 8304 1636 8356
rect 2688 8304 2740 8356
rect 8576 8304 8628 8356
rect 10692 8304 10744 8356
rect 2044 8279 2096 8288
rect 2044 8245 2053 8279
rect 2053 8245 2087 8279
rect 2087 8245 2096 8279
rect 2044 8236 2096 8245
rect 4528 8279 4580 8288
rect 4528 8245 4537 8279
rect 4537 8245 4571 8279
rect 4571 8245 4580 8279
rect 4528 8236 4580 8245
rect 9036 8236 9088 8288
rect 9496 8236 9548 8288
rect 9588 8236 9640 8288
rect 9956 8236 10008 8288
rect 2169 8134 2221 8186
rect 2233 8134 2285 8186
rect 2297 8134 2349 8186
rect 2361 8134 2413 8186
rect 2425 8134 2477 8186
rect 4607 8134 4659 8186
rect 4671 8134 4723 8186
rect 4735 8134 4787 8186
rect 4799 8134 4851 8186
rect 4863 8134 4915 8186
rect 7045 8134 7097 8186
rect 7109 8134 7161 8186
rect 7173 8134 7225 8186
rect 7237 8134 7289 8186
rect 7301 8134 7353 8186
rect 9483 8134 9535 8186
rect 9547 8134 9599 8186
rect 9611 8134 9663 8186
rect 9675 8134 9727 8186
rect 9739 8134 9791 8186
rect 2504 8032 2556 8084
rect 2964 8075 3016 8084
rect 2964 8041 2973 8075
rect 2973 8041 3007 8075
rect 3007 8041 3016 8075
rect 2964 8032 3016 8041
rect 1400 7964 1452 8016
rect 2136 7964 2188 8016
rect 3332 8032 3384 8084
rect 4252 8032 4304 8084
rect 6828 8032 6880 8084
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1860 7896 1912 7948
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 6460 7964 6512 8016
rect 6736 7964 6788 8016
rect 8024 7964 8076 8016
rect 2504 7828 2556 7880
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 3148 7828 3200 7880
rect 3240 7828 3292 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4528 7828 4580 7880
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 1584 7692 1636 7744
rect 2044 7692 2096 7744
rect 2964 7760 3016 7812
rect 3608 7803 3660 7812
rect 3608 7769 3617 7803
rect 3617 7769 3651 7803
rect 3651 7769 3660 7803
rect 3608 7760 3660 7769
rect 5632 7828 5684 7880
rect 5816 7828 5868 7880
rect 6460 7871 6512 7880
rect 6460 7837 6463 7871
rect 6463 7837 6512 7871
rect 6460 7828 6512 7837
rect 6552 7828 6604 7880
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 6184 7803 6236 7812
rect 6184 7769 6193 7803
rect 6193 7769 6227 7803
rect 6227 7769 6236 7803
rect 6184 7760 6236 7769
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 9036 7964 9088 8016
rect 9404 8032 9456 8084
rect 9864 8032 9916 8084
rect 10232 7964 10284 8016
rect 8392 7828 8444 7880
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 8852 7896 8904 7948
rect 8668 7760 8720 7812
rect 9496 7828 9548 7880
rect 9956 7828 10008 7880
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 4160 7692 4212 7744
rect 4436 7692 4488 7744
rect 6736 7692 6788 7744
rect 7104 7692 7156 7744
rect 8852 7692 8904 7744
rect 9220 7803 9272 7812
rect 9220 7769 9229 7803
rect 9229 7769 9263 7803
rect 9263 7769 9272 7803
rect 9220 7760 9272 7769
rect 9312 7803 9364 7812
rect 9312 7769 9321 7803
rect 9321 7769 9355 7803
rect 9355 7769 9364 7803
rect 9312 7760 9364 7769
rect 10048 7760 10100 7812
rect 9496 7692 9548 7744
rect 2829 7590 2881 7642
rect 2893 7590 2945 7642
rect 2957 7590 3009 7642
rect 3021 7590 3073 7642
rect 3085 7590 3137 7642
rect 5267 7590 5319 7642
rect 5331 7590 5383 7642
rect 5395 7590 5447 7642
rect 5459 7590 5511 7642
rect 5523 7590 5575 7642
rect 7705 7590 7757 7642
rect 7769 7590 7821 7642
rect 7833 7590 7885 7642
rect 7897 7590 7949 7642
rect 7961 7590 8013 7642
rect 10143 7590 10195 7642
rect 10207 7590 10259 7642
rect 10271 7590 10323 7642
rect 10335 7590 10387 7642
rect 10399 7590 10451 7642
rect 1676 7488 1728 7540
rect 2044 7488 2096 7540
rect 3240 7488 3292 7540
rect 3332 7488 3384 7540
rect 848 7352 900 7404
rect 1584 7352 1636 7404
rect 2596 7463 2648 7472
rect 2596 7429 2605 7463
rect 2605 7429 2639 7463
rect 2639 7429 2648 7463
rect 2596 7420 2648 7429
rect 2688 7420 2740 7472
rect 3792 7420 3844 7472
rect 4252 7488 4304 7540
rect 5172 7488 5224 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 3332 7352 3384 7404
rect 3608 7352 3660 7404
rect 4988 7420 5040 7472
rect 7380 7488 7432 7540
rect 8668 7488 8720 7540
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 6736 7395 6788 7404
rect 6736 7361 6742 7395
rect 6742 7361 6776 7395
rect 6776 7361 6788 7395
rect 6736 7352 6788 7361
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 8852 7463 8904 7472
rect 8852 7429 8861 7463
rect 8861 7429 8895 7463
rect 8895 7429 8904 7463
rect 8852 7420 8904 7429
rect 9496 7488 9548 7540
rect 8392 7352 8444 7404
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 6184 7284 6236 7336
rect 7012 7284 7064 7336
rect 9036 7352 9088 7404
rect 9220 7352 9272 7404
rect 9864 7420 9916 7472
rect 10232 7352 10284 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 4528 7216 4580 7268
rect 6460 7216 6512 7268
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 9128 7216 9180 7268
rect 4252 7148 4304 7200
rect 2169 7046 2221 7098
rect 2233 7046 2285 7098
rect 2297 7046 2349 7098
rect 2361 7046 2413 7098
rect 2425 7046 2477 7098
rect 4607 7046 4659 7098
rect 4671 7046 4723 7098
rect 4735 7046 4787 7098
rect 4799 7046 4851 7098
rect 4863 7046 4915 7098
rect 7045 7046 7097 7098
rect 7109 7046 7161 7098
rect 7173 7046 7225 7098
rect 7237 7046 7289 7098
rect 7301 7046 7353 7098
rect 9483 7046 9535 7098
rect 9547 7046 9599 7098
rect 9611 7046 9663 7098
rect 9675 7046 9727 7098
rect 9739 7046 9791 7098
rect 1952 6944 2004 6996
rect 5816 6944 5868 6996
rect 8576 6944 8628 6996
rect 6000 6876 6052 6928
rect 1860 6808 1912 6860
rect 2228 6808 2280 6860
rect 1768 6672 1820 6724
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 9864 6876 9916 6928
rect 8852 6808 8904 6860
rect 10048 6808 10100 6860
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 6184 6672 6236 6724
rect 7380 6672 7432 6724
rect 9956 6740 10008 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 9220 6604 9272 6656
rect 2829 6502 2881 6554
rect 2893 6502 2945 6554
rect 2957 6502 3009 6554
rect 3021 6502 3073 6554
rect 3085 6502 3137 6554
rect 5267 6502 5319 6554
rect 5331 6502 5383 6554
rect 5395 6502 5447 6554
rect 5459 6502 5511 6554
rect 5523 6502 5575 6554
rect 7705 6502 7757 6554
rect 7769 6502 7821 6554
rect 7833 6502 7885 6554
rect 7897 6502 7949 6554
rect 7961 6502 8013 6554
rect 10143 6502 10195 6554
rect 10207 6502 10259 6554
rect 10271 6502 10323 6554
rect 10335 6502 10387 6554
rect 10399 6502 10451 6554
rect 2228 6375 2280 6384
rect 2228 6341 2237 6375
rect 2237 6341 2271 6375
rect 2271 6341 2280 6375
rect 2228 6332 2280 6341
rect 2780 6400 2832 6452
rect 3608 6400 3660 6452
rect 9128 6400 9180 6452
rect 4160 6375 4212 6384
rect 4160 6341 4169 6375
rect 4169 6341 4203 6375
rect 4203 6341 4212 6375
rect 4160 6332 4212 6341
rect 6736 6332 6788 6384
rect 848 6264 900 6316
rect 3056 6264 3108 6316
rect 3700 6264 3752 6316
rect 8760 6264 8812 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 10416 6307 10468 6316
rect 10416 6273 10425 6307
rect 10425 6273 10459 6307
rect 10459 6273 10468 6307
rect 10416 6264 10468 6273
rect 5080 6196 5132 6248
rect 8392 6196 8444 6248
rect 10048 6196 10100 6248
rect 3424 6128 3476 6180
rect 9404 6128 9456 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 4436 6060 4488 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 4988 6060 5040 6112
rect 5448 6103 5500 6112
rect 5448 6069 5457 6103
rect 5457 6069 5491 6103
rect 5491 6069 5500 6103
rect 5448 6060 5500 6069
rect 2169 5958 2221 6010
rect 2233 5958 2285 6010
rect 2297 5958 2349 6010
rect 2361 5958 2413 6010
rect 2425 5958 2477 6010
rect 4607 5958 4659 6010
rect 4671 5958 4723 6010
rect 4735 5958 4787 6010
rect 4799 5958 4851 6010
rect 4863 5958 4915 6010
rect 7045 5958 7097 6010
rect 7109 5958 7161 6010
rect 7173 5958 7225 6010
rect 7237 5958 7289 6010
rect 7301 5958 7353 6010
rect 9483 5958 9535 6010
rect 9547 5958 9599 6010
rect 9611 5958 9663 6010
rect 9675 5958 9727 6010
rect 9739 5958 9791 6010
rect 1952 5788 2004 5840
rect 2044 5763 2096 5772
rect 2044 5729 2053 5763
rect 2053 5729 2087 5763
rect 2087 5729 2096 5763
rect 2044 5720 2096 5729
rect 2596 5720 2648 5772
rect 3148 5788 3200 5840
rect 2964 5720 3016 5772
rect 3240 5720 3292 5772
rect 5172 5856 5224 5908
rect 6552 5856 6604 5908
rect 7288 5856 7340 5908
rect 7656 5856 7708 5908
rect 8576 5856 8628 5908
rect 8944 5856 8996 5908
rect 3792 5788 3844 5840
rect 1676 5627 1728 5636
rect 1676 5593 1685 5627
rect 1685 5593 1719 5627
rect 1719 5593 1728 5627
rect 1676 5584 1728 5593
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 1400 5559 1452 5568
rect 1400 5525 1409 5559
rect 1409 5525 1443 5559
rect 1443 5525 1452 5559
rect 1400 5516 1452 5525
rect 3332 5652 3384 5704
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 4160 5720 4212 5772
rect 5724 5788 5776 5840
rect 5908 5788 5960 5840
rect 6920 5788 6972 5840
rect 9956 5831 10008 5840
rect 9956 5797 9965 5831
rect 9965 5797 9999 5831
rect 9999 5797 10008 5831
rect 9956 5788 10008 5797
rect 4988 5720 5040 5772
rect 2688 5584 2740 5636
rect 2780 5584 2832 5636
rect 3056 5584 3108 5636
rect 4528 5652 4580 5704
rect 5632 5720 5684 5772
rect 6644 5720 6696 5772
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 3148 5516 3200 5568
rect 3792 5516 3844 5568
rect 4436 5516 4488 5568
rect 5632 5516 5684 5568
rect 6460 5516 6512 5568
rect 7472 5584 7524 5636
rect 8852 5652 8904 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9404 5652 9456 5704
rect 8024 5584 8076 5636
rect 7564 5516 7616 5568
rect 8208 5516 8260 5568
rect 8576 5627 8628 5636
rect 8576 5593 8585 5627
rect 8585 5593 8619 5627
rect 8619 5593 8628 5627
rect 8576 5584 8628 5593
rect 10600 5652 10652 5704
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 2829 5414 2881 5466
rect 2893 5414 2945 5466
rect 2957 5414 3009 5466
rect 3021 5414 3073 5466
rect 3085 5414 3137 5466
rect 5267 5414 5319 5466
rect 5331 5414 5383 5466
rect 5395 5414 5447 5466
rect 5459 5414 5511 5466
rect 5523 5414 5575 5466
rect 7705 5414 7757 5466
rect 7769 5414 7821 5466
rect 7833 5414 7885 5466
rect 7897 5414 7949 5466
rect 7961 5414 8013 5466
rect 10143 5414 10195 5466
rect 10207 5414 10259 5466
rect 10271 5414 10323 5466
rect 10335 5414 10387 5466
rect 10399 5414 10451 5466
rect 1308 5312 1360 5364
rect 1676 5312 1728 5364
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 1400 5244 1452 5296
rect 5172 5312 5224 5364
rect 7196 5312 7248 5364
rect 7472 5355 7524 5364
rect 7472 5321 7481 5355
rect 7481 5321 7515 5355
rect 7515 5321 7524 5355
rect 7472 5312 7524 5321
rect 3240 5176 3292 5228
rect 3424 5176 3476 5228
rect 4160 5244 4212 5296
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 2504 5108 2556 5160
rect 6460 5219 6512 5228
rect 6460 5185 6469 5219
rect 6469 5185 6503 5219
rect 6503 5185 6512 5219
rect 6460 5176 6512 5185
rect 8208 5244 8260 5296
rect 7472 5176 7524 5228
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 8392 5176 8444 5228
rect 8576 5176 8628 5228
rect 9312 5176 9364 5228
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 4436 5108 4488 5160
rect 6736 5108 6788 5160
rect 3240 5040 3292 5092
rect 3332 4972 3384 5024
rect 8760 5040 8812 5092
rect 8852 5040 8904 5092
rect 9312 5083 9364 5092
rect 9312 5049 9321 5083
rect 9321 5049 9355 5083
rect 9355 5049 9364 5083
rect 9312 5040 9364 5049
rect 6920 4972 6972 5024
rect 7288 4972 7340 5024
rect 7656 4972 7708 5024
rect 2169 4870 2221 4922
rect 2233 4870 2285 4922
rect 2297 4870 2349 4922
rect 2361 4870 2413 4922
rect 2425 4870 2477 4922
rect 4607 4870 4659 4922
rect 4671 4870 4723 4922
rect 4735 4870 4787 4922
rect 4799 4870 4851 4922
rect 4863 4870 4915 4922
rect 7045 4870 7097 4922
rect 7109 4870 7161 4922
rect 7173 4870 7225 4922
rect 7237 4870 7289 4922
rect 7301 4870 7353 4922
rect 9483 4870 9535 4922
rect 9547 4870 9599 4922
rect 9611 4870 9663 4922
rect 9675 4870 9727 4922
rect 9739 4870 9791 4922
rect 2504 4768 2556 4820
rect 5816 4768 5868 4820
rect 6736 4768 6788 4820
rect 7564 4768 7616 4820
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 7380 4632 7432 4684
rect 848 4564 900 4616
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 6828 4564 6880 4616
rect 8024 4564 8076 4616
rect 8300 4632 8352 4684
rect 8944 4632 8996 4684
rect 9312 4632 9364 4684
rect 8300 4496 8352 4548
rect 8208 4428 8260 4480
rect 9036 4564 9088 4616
rect 2829 4326 2881 4378
rect 2893 4326 2945 4378
rect 2957 4326 3009 4378
rect 3021 4326 3073 4378
rect 3085 4326 3137 4378
rect 5267 4326 5319 4378
rect 5331 4326 5383 4378
rect 5395 4326 5447 4378
rect 5459 4326 5511 4378
rect 5523 4326 5575 4378
rect 7705 4326 7757 4378
rect 7769 4326 7821 4378
rect 7833 4326 7885 4378
rect 7897 4326 7949 4378
rect 7961 4326 8013 4378
rect 10143 4326 10195 4378
rect 10207 4326 10259 4378
rect 10271 4326 10323 4378
rect 10335 4326 10387 4378
rect 10399 4326 10451 4378
rect 4344 4088 4396 4140
rect 5724 4199 5776 4208
rect 5724 4165 5733 4199
rect 5733 4165 5767 4199
rect 5767 4165 5776 4199
rect 5724 4156 5776 4165
rect 6736 4156 6788 4208
rect 7380 4156 7432 4208
rect 5080 4020 5132 4072
rect 4436 3952 4488 4004
rect 5632 4020 5684 4072
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 9864 4088 9916 4140
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 8852 4020 8904 4072
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 4528 3884 4580 3936
rect 4988 3884 5040 3936
rect 5632 3884 5684 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 9404 3884 9456 3936
rect 2169 3782 2221 3834
rect 2233 3782 2285 3834
rect 2297 3782 2349 3834
rect 2361 3782 2413 3834
rect 2425 3782 2477 3834
rect 4607 3782 4659 3834
rect 4671 3782 4723 3834
rect 4735 3782 4787 3834
rect 4799 3782 4851 3834
rect 4863 3782 4915 3834
rect 7045 3782 7097 3834
rect 7109 3782 7161 3834
rect 7173 3782 7225 3834
rect 7237 3782 7289 3834
rect 7301 3782 7353 3834
rect 9483 3782 9535 3834
rect 9547 3782 9599 3834
rect 9611 3782 9663 3834
rect 9675 3782 9727 3834
rect 9739 3782 9791 3834
rect 2688 3680 2740 3732
rect 4620 3680 4672 3732
rect 2780 3612 2832 3664
rect 848 3544 900 3596
rect 1768 3544 1820 3596
rect 4528 3612 4580 3664
rect 6644 3680 6696 3732
rect 9128 3680 9180 3732
rect 10048 3680 10100 3732
rect 8392 3612 8444 3664
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 3516 3544 3568 3553
rect 4160 3544 4212 3596
rect 3332 3476 3384 3528
rect 4620 3544 4672 3596
rect 5172 3544 5224 3596
rect 7380 3544 7432 3596
rect 3424 3408 3476 3460
rect 4528 3476 4580 3528
rect 4988 3476 5040 3528
rect 5080 3476 5132 3528
rect 5724 3476 5776 3528
rect 7564 3476 7616 3528
rect 8852 3544 8904 3596
rect 2228 3340 2280 3392
rect 3240 3340 3292 3392
rect 6644 3408 6696 3460
rect 4436 3340 4488 3392
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 7564 3340 7616 3392
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 9404 3408 9456 3460
rect 8944 3340 8996 3392
rect 2829 3238 2881 3290
rect 2893 3238 2945 3290
rect 2957 3238 3009 3290
rect 3021 3238 3073 3290
rect 3085 3238 3137 3290
rect 5267 3238 5319 3290
rect 5331 3238 5383 3290
rect 5395 3238 5447 3290
rect 5459 3238 5511 3290
rect 5523 3238 5575 3290
rect 7705 3238 7757 3290
rect 7769 3238 7821 3290
rect 7833 3238 7885 3290
rect 7897 3238 7949 3290
rect 7961 3238 8013 3290
rect 10143 3238 10195 3290
rect 10207 3238 10259 3290
rect 10271 3238 10323 3290
rect 10335 3238 10387 3290
rect 10399 3238 10451 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 2780 3136 2832 3145
rect 3424 3136 3476 3188
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 3240 3068 3292 3120
rect 4344 3068 4396 3120
rect 5080 3136 5132 3188
rect 5172 3136 5224 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7380 3136 7432 3188
rect 8944 3136 8996 3188
rect 9312 3136 9364 3188
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 4068 3000 4120 3052
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 4160 2932 4212 2984
rect 3332 2864 3384 2916
rect 4344 2864 4396 2916
rect 5816 3068 5868 3120
rect 7472 3068 7524 3120
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 8668 3068 8720 3120
rect 9588 3136 9640 3188
rect 9680 3136 9732 3188
rect 8484 3000 8536 3052
rect 8392 2975 8444 2984
rect 8392 2941 8401 2975
rect 8401 2941 8435 2975
rect 8435 2941 8444 2975
rect 9496 3068 9548 3120
rect 9956 3068 10008 3120
rect 9404 3000 9456 3052
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 9864 3000 9916 3052
rect 8392 2932 8444 2941
rect 9496 2932 9548 2984
rect 9220 2864 9272 2916
rect 5632 2796 5684 2848
rect 7840 2796 7892 2848
rect 8484 2796 8536 2848
rect 2169 2694 2221 2746
rect 2233 2694 2285 2746
rect 2297 2694 2349 2746
rect 2361 2694 2413 2746
rect 2425 2694 2477 2746
rect 4607 2694 4659 2746
rect 4671 2694 4723 2746
rect 4735 2694 4787 2746
rect 4799 2694 4851 2746
rect 4863 2694 4915 2746
rect 7045 2694 7097 2746
rect 7109 2694 7161 2746
rect 7173 2694 7225 2746
rect 7237 2694 7289 2746
rect 7301 2694 7353 2746
rect 9483 2694 9535 2746
rect 9547 2694 9599 2746
rect 9611 2694 9663 2746
rect 9675 2694 9727 2746
rect 9739 2694 9791 2746
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 4436 2592 4488 2644
rect 6460 2592 6512 2644
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 9220 2592 9272 2644
rect 9312 2635 9364 2644
rect 9312 2601 9321 2635
rect 9321 2601 9355 2635
rect 9355 2601 9364 2635
rect 9312 2592 9364 2601
rect 9864 2592 9916 2644
rect 3884 2388 3936 2440
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 5724 2388 5776 2440
rect 6460 2388 6512 2440
rect 6920 2388 6972 2440
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8392 2388 8444 2440
rect 9036 2388 9088 2440
rect 9680 2388 9732 2440
rect 5172 2320 5224 2372
rect 7104 2252 7156 2304
rect 7564 2252 7616 2304
rect 2829 2150 2881 2202
rect 2893 2150 2945 2202
rect 2957 2150 3009 2202
rect 3021 2150 3073 2202
rect 3085 2150 3137 2202
rect 5267 2150 5319 2202
rect 5331 2150 5383 2202
rect 5395 2150 5447 2202
rect 5459 2150 5511 2202
rect 5523 2150 5575 2202
rect 7705 2150 7757 2202
rect 7769 2150 7821 2202
rect 7833 2150 7885 2202
rect 7897 2150 7949 2202
rect 7961 2150 8013 2202
rect 10143 2150 10195 2202
rect 10207 2150 10259 2202
rect 10271 2150 10323 2202
rect 10335 2150 10387 2202
rect 10399 2150 10451 2202
<< metal2 >>
rect 3882 13342 3938 14142
rect 4526 13342 4582 14142
rect 5814 13342 5870 14142
rect 7102 13342 7158 14142
rect 7746 13342 7802 14142
rect 7852 13382 8156 13410
rect 2169 11452 2477 11461
rect 2169 11450 2175 11452
rect 2231 11450 2255 11452
rect 2311 11450 2335 11452
rect 2391 11450 2415 11452
rect 2471 11450 2477 11452
rect 2231 11398 2233 11450
rect 2413 11398 2415 11450
rect 2169 11396 2175 11398
rect 2231 11396 2255 11398
rect 2311 11396 2335 11398
rect 2391 11396 2415 11398
rect 2471 11396 2477 11398
rect 2169 11387 2477 11396
rect 3896 11150 3924 13342
rect 4540 11218 4568 13342
rect 4607 11452 4915 11461
rect 4607 11450 4613 11452
rect 4669 11450 4693 11452
rect 4749 11450 4773 11452
rect 4829 11450 4853 11452
rect 4909 11450 4915 11452
rect 4669 11398 4671 11450
rect 4851 11398 4853 11450
rect 4607 11396 4613 11398
rect 4669 11396 4693 11398
rect 4749 11396 4773 11398
rect 4829 11396 4853 11398
rect 4909 11396 4915 11398
rect 4607 11387 4915 11396
rect 5828 11354 5856 13342
rect 7116 11898 7144 13342
rect 7760 13274 7788 13342
rect 7852 13274 7880 13382
rect 7760 13246 7880 13274
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7045 11452 7353 11461
rect 7045 11450 7051 11452
rect 7107 11450 7131 11452
rect 7187 11450 7211 11452
rect 7267 11450 7291 11452
rect 7347 11450 7353 11452
rect 7107 11398 7109 11450
rect 7289 11398 7291 11450
rect 7045 11396 7051 11398
rect 7107 11396 7131 11398
rect 7187 11396 7211 11398
rect 7267 11396 7291 11398
rect 7347 11396 7353 11398
rect 7045 11387 7353 11396
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 2829 10908 3137 10917
rect 2829 10906 2835 10908
rect 2891 10906 2915 10908
rect 2971 10906 2995 10908
rect 3051 10906 3075 10908
rect 3131 10906 3137 10908
rect 2891 10854 2893 10906
rect 3073 10854 3075 10906
rect 2829 10852 2835 10854
rect 2891 10852 2915 10854
rect 2971 10852 2995 10854
rect 3051 10852 3075 10854
rect 3131 10852 3137 10854
rect 2829 10843 3137 10852
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 1676 10464 1728 10470
rect 900 10432 902 10441
rect 1676 10406 1728 10412
rect 846 10367 902 10376
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 846 9072 902 9081
rect 846 9007 902 9016
rect 860 8974 888 9007
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 1412 8022 1440 10066
rect 1688 10062 1716 10406
rect 2056 10266 2084 10610
rect 2169 10364 2477 10373
rect 2169 10362 2175 10364
rect 2231 10362 2255 10364
rect 2311 10362 2335 10364
rect 2391 10362 2415 10364
rect 2471 10362 2477 10364
rect 2231 10310 2233 10362
rect 2413 10310 2415 10362
rect 2169 10308 2175 10310
rect 2231 10308 2255 10310
rect 2311 10308 2335 10310
rect 2391 10308 2415 10310
rect 2471 10308 2477 10310
rect 2169 10299 2477 10308
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2792 10198 2820 10610
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1780 9450 1808 9930
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1400 8016 1452 8022
rect 1400 7958 1452 7964
rect 1596 7886 1624 8298
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 846 7440 902 7449
rect 1596 7410 1624 7686
rect 1688 7546 1716 8434
rect 1872 7954 1900 9930
rect 2148 9722 2176 9998
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2516 9654 2544 9998
rect 2792 9908 2820 10134
rect 2700 9880 2820 9908
rect 2700 9704 2728 9880
rect 2829 9820 3137 9829
rect 2829 9818 2835 9820
rect 2891 9818 2915 9820
rect 2971 9818 2995 9820
rect 3051 9818 3075 9820
rect 3131 9818 3137 9820
rect 2891 9766 2893 9818
rect 3073 9766 3075 9818
rect 2829 9764 2835 9766
rect 2891 9764 2915 9766
rect 2971 9764 2995 9766
rect 3051 9764 3075 9766
rect 3131 9764 3137 9766
rect 2829 9755 3137 9764
rect 2700 9676 2820 9704
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1964 8498 1992 9522
rect 2792 9382 2820 9676
rect 3252 9586 3280 10406
rect 3436 10062 3464 10678
rect 3896 10606 3924 10950
rect 4264 10674 4292 10950
rect 5092 10810 5120 10950
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5184 10690 5212 11086
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 5267 10908 5575 10917
rect 5267 10906 5273 10908
rect 5329 10906 5353 10908
rect 5409 10906 5433 10908
rect 5489 10906 5513 10908
rect 5569 10906 5575 10908
rect 5329 10854 5331 10906
rect 5511 10854 5513 10906
rect 5267 10852 5273 10854
rect 5329 10852 5353 10854
rect 5409 10852 5433 10854
rect 5489 10852 5513 10854
rect 5569 10852 5575 10854
rect 5267 10843 5575 10852
rect 6472 10810 6500 11018
rect 7116 10810 7144 11154
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7392 10742 7420 11086
rect 7484 10810 7512 11086
rect 7705 10908 8013 10917
rect 7705 10906 7711 10908
rect 7767 10906 7791 10908
rect 7847 10906 7871 10908
rect 7927 10906 7951 10908
rect 8007 10906 8013 10908
rect 7767 10854 7769 10906
rect 7949 10854 7951 10906
rect 7705 10852 7711 10854
rect 7767 10852 7791 10854
rect 7847 10852 7871 10854
rect 7927 10852 7951 10854
rect 8007 10852 8013 10854
rect 7705 10843 8013 10852
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 5264 10736 5316 10742
rect 5184 10684 5264 10690
rect 5184 10678 5316 10684
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 4252 10668 4304 10674
rect 5184 10662 5304 10678
rect 4252 10610 4304 10616
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3344 9382 3372 9930
rect 3436 9586 3464 9998
rect 3804 9654 3832 10202
rect 3896 10062 3924 10542
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4080 10198 4108 10474
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3896 9586 3924 9998
rect 4172 9586 4200 10066
rect 4448 10062 4476 10406
rect 4607 10364 4915 10373
rect 4607 10362 4613 10364
rect 4669 10362 4693 10364
rect 4749 10362 4773 10364
rect 4829 10362 4853 10364
rect 4909 10362 4915 10364
rect 4669 10310 4671 10362
rect 4851 10310 4853 10362
rect 4607 10308 4613 10310
rect 4669 10308 4693 10310
rect 4749 10308 4773 10310
rect 4829 10308 4853 10310
rect 4909 10308 4915 10310
rect 4607 10299 4915 10308
rect 5276 10198 5304 10662
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10198 5396 10406
rect 5552 10266 5580 10610
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5828 10130 5856 10406
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 6196 10062 6224 10406
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 2169 9276 2477 9285
rect 2169 9274 2175 9276
rect 2231 9274 2255 9276
rect 2311 9274 2335 9276
rect 2391 9274 2415 9276
rect 2471 9274 2477 9276
rect 2231 9222 2233 9274
rect 2413 9222 2415 9274
rect 2169 9220 2175 9222
rect 2231 9220 2255 9222
rect 2311 9220 2335 9222
rect 2391 9220 2415 9222
rect 2471 9220 2477 9222
rect 2169 9211 2477 9220
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 2829 8732 3137 8741
rect 2829 8730 2835 8732
rect 2891 8730 2915 8732
rect 2971 8730 2995 8732
rect 3051 8730 3075 8732
rect 3131 8730 3137 8732
rect 2891 8678 2893 8730
rect 3073 8678 3075 8730
rect 2829 8676 2835 8678
rect 2891 8676 2915 8678
rect 2971 8676 2995 8678
rect 3051 8676 3075 8678
rect 3131 8676 3137 8678
rect 2829 8667 3137 8676
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 1860 7948 1912 7954
rect 1780 7908 1860 7936
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 846 7375 848 7384
rect 900 7375 902 7384
rect 1584 7404 1636 7410
rect 848 7346 900 7352
rect 1584 7346 1636 7352
rect 1780 6730 1808 7908
rect 1860 7890 1912 7896
rect 1964 7834 1992 8434
rect 2424 8378 2452 8434
rect 2424 8350 2544 8378
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2056 7954 2084 8230
rect 2169 8188 2477 8197
rect 2169 8186 2175 8188
rect 2231 8186 2255 8188
rect 2311 8186 2335 8188
rect 2391 8186 2415 8188
rect 2471 8186 2477 8188
rect 2231 8134 2233 8186
rect 2413 8134 2415 8186
rect 2169 8132 2175 8134
rect 2231 8132 2255 8134
rect 2311 8132 2335 8134
rect 2391 8132 2415 8134
rect 2471 8132 2477 8134
rect 2169 8123 2477 8132
rect 2516 8090 2544 8350
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 1872 7806 1992 7834
rect 1872 6866 1900 7806
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2056 7546 2084 7686
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2148 7426 2176 7958
rect 2516 7886 2544 8026
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2608 7478 2636 8434
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 7834 2728 8298
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7880 2924 7886
rect 2700 7828 2872 7834
rect 2700 7822 2924 7828
rect 2700 7806 2912 7822
rect 2976 7818 3004 8026
rect 3252 7970 3280 8774
rect 3344 8090 3372 9318
rect 4264 8090 4292 9862
rect 4632 9722 4660 9998
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4816 9654 4844 9862
rect 5267 9820 5575 9829
rect 5267 9818 5273 9820
rect 5329 9818 5353 9820
rect 5409 9818 5433 9820
rect 5489 9818 5513 9820
rect 5569 9818 5575 9820
rect 5329 9766 5331 9818
rect 5511 9766 5513 9818
rect 5267 9764 5273 9766
rect 5329 9764 5353 9766
rect 5409 9764 5433 9766
rect 5489 9764 5513 9766
rect 5569 9764 5575 9766
rect 5267 9755 5575 9764
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4607 9276 4915 9285
rect 4607 9274 4613 9276
rect 4669 9274 4693 9276
rect 4749 9274 4773 9276
rect 4829 9274 4853 9276
rect 4909 9274 4915 9276
rect 4669 9222 4671 9274
rect 4851 9222 4853 9274
rect 4607 9220 4613 9222
rect 4669 9220 4693 9222
rect 4749 9220 4773 9222
rect 4829 9220 4853 9222
rect 4909 9220 4915 9222
rect 4607 9211 4915 9220
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3160 7942 3372 7970
rect 3160 7886 3188 7942
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2964 7812 3016 7818
rect 2700 7478 2728 7806
rect 2964 7754 3016 7760
rect 2829 7644 3137 7653
rect 2829 7642 2835 7644
rect 2891 7642 2915 7644
rect 2971 7642 2995 7644
rect 3051 7642 3075 7644
rect 3131 7642 3137 7644
rect 2891 7590 2893 7642
rect 3073 7590 3075 7642
rect 2829 7588 2835 7590
rect 2891 7588 2915 7590
rect 2971 7588 2995 7590
rect 3051 7588 3075 7590
rect 3131 7588 3137 7590
rect 2829 7579 3137 7588
rect 3252 7546 3280 7822
rect 3344 7546 3372 7942
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 1964 7398 2176 7426
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 3344 7410 3372 7482
rect 3620 7410 3648 7754
rect 3804 7478 3832 7822
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3332 7404 3384 7410
rect 1964 7002 1992 7398
rect 3332 7346 3384 7352
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 2169 7100 2477 7109
rect 2169 7098 2175 7100
rect 2231 7098 2255 7100
rect 2311 7098 2335 7100
rect 2391 7098 2415 7100
rect 2471 7098 2477 7100
rect 2231 7046 2233 7098
rect 2413 7046 2415 7098
rect 2169 7044 2175 7046
rect 2231 7044 2255 7046
rect 2311 7044 2335 7046
rect 2391 7044 2415 7046
rect 2471 7044 2477 7046
rect 2169 7035 2477 7044
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1780 5642 1808 6666
rect 1964 5846 1992 6938
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2240 6390 2268 6802
rect 2829 6556 3137 6565
rect 2829 6554 2835 6556
rect 2891 6554 2915 6556
rect 2971 6554 2995 6556
rect 3051 6554 3075 6556
rect 3131 6554 3137 6556
rect 2891 6502 2893 6554
rect 3073 6502 3075 6554
rect 2829 6500 2835 6502
rect 2891 6500 2915 6502
rect 2971 6500 2995 6502
rect 3051 6500 3075 6502
rect 3131 6500 3137 6502
rect 2829 6491 3137 6500
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 2056 5778 2084 6054
rect 2169 6012 2477 6021
rect 2169 6010 2175 6012
rect 2231 6010 2255 6012
rect 2311 6010 2335 6012
rect 2391 6010 2415 6012
rect 2471 6010 2477 6012
rect 2231 5958 2233 6010
rect 2413 5958 2415 6010
rect 2169 5956 2175 5958
rect 2231 5956 2255 5958
rect 2311 5956 2335 5958
rect 2391 5956 2415 5958
rect 2471 5956 2477 5958
rect 2169 5947 2477 5956
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1400 5568 1452 5574
rect 1306 5536 1362 5545
rect 1400 5510 1452 5516
rect 1306 5471 1362 5480
rect 1320 5370 1348 5471
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1412 5302 1440 5510
rect 1688 5370 1716 5578
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1400 5296 1452 5302
rect 1400 5238 1452 5244
rect 846 4720 902 4729
rect 846 4655 902 4664
rect 860 4622 888 4655
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 846 3632 902 3641
rect 1780 3602 1808 5578
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2169 4924 2477 4933
rect 2169 4922 2175 4924
rect 2231 4922 2255 4924
rect 2311 4922 2335 4924
rect 2391 4922 2415 4924
rect 2471 4922 2477 4924
rect 2231 4870 2233 4922
rect 2413 4870 2415 4922
rect 2169 4868 2175 4870
rect 2231 4868 2255 4870
rect 2311 4868 2335 4870
rect 2391 4868 2415 4870
rect 2471 4868 2477 4870
rect 2169 4859 2477 4868
rect 2516 4826 2544 5102
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2169 3836 2477 3845
rect 2169 3834 2175 3836
rect 2231 3834 2255 3836
rect 2311 3834 2335 3836
rect 2391 3834 2415 3836
rect 2471 3834 2477 3836
rect 2231 3782 2233 3834
rect 2413 3782 2415 3834
rect 2169 3780 2175 3782
rect 2231 3780 2255 3782
rect 2311 3780 2335 3782
rect 2391 3780 2415 3782
rect 2471 3780 2477 3782
rect 2169 3771 2477 3780
rect 2608 3641 2636 5714
rect 2792 5642 2820 6394
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2964 5772 3016 5778
rect 3068 5760 3096 6258
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3016 5732 3096 5760
rect 2964 5714 3016 5720
rect 3068 5642 3096 5732
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2700 4162 2728 5578
rect 3160 5574 3188 5782
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2829 5468 3137 5477
rect 2829 5466 2835 5468
rect 2891 5466 2915 5468
rect 2971 5466 2995 5468
rect 3051 5466 3075 5468
rect 3131 5466 3137 5468
rect 2891 5414 2893 5466
rect 3073 5414 3075 5466
rect 2829 5412 2835 5414
rect 2891 5412 2915 5414
rect 2971 5412 2995 5414
rect 3051 5412 3075 5414
rect 3131 5412 3137 5414
rect 2829 5403 3137 5412
rect 3252 5234 3280 5714
rect 3436 5710 3464 6122
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 5098 3280 5170
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3344 5030 3372 5646
rect 3436 5234 3464 5646
rect 3620 5370 3648 6394
rect 4172 6390 4200 7686
rect 4264 7546 4292 8026
rect 4540 7886 4568 8230
rect 4607 8188 4915 8197
rect 4607 8186 4613 8188
rect 4669 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4915 8188
rect 4669 8134 4671 8186
rect 4851 8134 4853 8186
rect 4607 8132 4613 8134
rect 4669 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4915 8134
rect 4607 8123 4915 8132
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4264 7206 4292 7482
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3712 5234 3740 6258
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3804 5574 3832 5782
rect 4172 5778 4200 6326
rect 4448 6118 4476 7686
rect 4540 7274 4568 7822
rect 4632 7290 4660 7890
rect 5000 7478 5028 9386
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 5092 7290 5120 9454
rect 5644 9042 5672 9658
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5267 8732 5575 8741
rect 5267 8730 5273 8732
rect 5329 8730 5353 8732
rect 5409 8730 5433 8732
rect 5489 8730 5513 8732
rect 5569 8730 5575 8732
rect 5329 8678 5331 8730
rect 5511 8678 5513 8730
rect 5267 8676 5273 8678
rect 5329 8676 5353 8678
rect 5409 8676 5433 8678
rect 5489 8676 5513 8678
rect 5569 8676 5575 8678
rect 5267 8667 5575 8676
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5184 7886 5212 8434
rect 5644 7886 5672 8978
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5184 7546 5212 7822
rect 5267 7644 5575 7653
rect 5267 7642 5273 7644
rect 5329 7642 5353 7644
rect 5409 7642 5433 7644
rect 5489 7642 5513 7644
rect 5569 7642 5575 7644
rect 5329 7590 5331 7642
rect 5511 7590 5513 7642
rect 5267 7588 5273 7590
rect 5329 7588 5353 7590
rect 5409 7588 5433 7590
rect 5489 7588 5513 7590
rect 5569 7588 5575 7590
rect 5267 7579 5575 7588
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4528 7268 4580 7274
rect 4632 7262 5120 7290
rect 4528 7210 4580 7216
rect 4607 7100 4915 7109
rect 4607 7098 4613 7100
rect 4669 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4915 7100
rect 4669 7046 4671 7098
rect 4851 7046 4853 7098
rect 4607 7044 4613 7046
rect 4669 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4915 7046
rect 4607 7035 4915 7044
rect 5092 6254 5120 7262
rect 5267 6556 5575 6565
rect 5267 6554 5273 6556
rect 5329 6554 5353 6556
rect 5409 6554 5433 6556
rect 5489 6554 5513 6556
rect 5569 6554 5575 6556
rect 5329 6502 5331 6554
rect 5511 6502 5513 6554
rect 5267 6500 5273 6502
rect 5329 6500 5353 6502
rect 5409 6500 5433 6502
rect 5489 6500 5513 6502
rect 5569 6500 5575 6502
rect 5267 6491 5575 6500
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 4172 5302 4200 5714
rect 4448 5574 4476 6054
rect 4540 5710 4568 6054
rect 4607 6012 4915 6021
rect 4607 6010 4613 6012
rect 4669 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4915 6012
rect 4669 5958 4671 6010
rect 4851 5958 4853 6010
rect 4607 5956 4613 5958
rect 4669 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4915 5958
rect 4607 5947 4915 5956
rect 5000 5778 5028 6054
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 4448 5166 4476 5510
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 4607 4924 4915 4933
rect 4607 4922 4613 4924
rect 4669 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4915 4924
rect 4669 4870 4671 4922
rect 4851 4870 4853 4922
rect 4607 4868 4613 4870
rect 4669 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4915 4870
rect 4607 4859 4915 4868
rect 2829 4380 3137 4389
rect 2829 4378 2835 4380
rect 2891 4378 2915 4380
rect 2971 4378 2995 4380
rect 3051 4378 3075 4380
rect 3131 4378 3137 4380
rect 2891 4326 2893 4378
rect 3073 4326 3075 4378
rect 2829 4324 2835 4326
rect 2891 4324 2915 4326
rect 2971 4324 2995 4326
rect 3051 4324 3075 4326
rect 3131 4324 3137 4326
rect 2829 4315 3137 4324
rect 2700 4134 2820 4162
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2594 3632 2650 3641
rect 846 3567 848 3576
rect 900 3567 902 3576
rect 1768 3596 1820 3602
rect 848 3538 900 3544
rect 2594 3567 2650 3576
rect 1768 3538 1820 3544
rect 2700 3534 2728 3674
rect 2792 3670 2820 4134
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4356 4026 4384 4082
rect 5092 4078 5120 6190
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5184 5658 5212 5850
rect 5460 5710 5488 6054
rect 5644 5778 5672 7822
rect 5828 7410 5856 7822
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 7002 5856 7346
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5264 5704 5316 5710
rect 5184 5652 5264 5658
rect 5184 5646 5316 5652
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5184 5630 5304 5646
rect 5184 5370 5212 5630
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5267 5468 5575 5477
rect 5267 5466 5273 5468
rect 5329 5466 5353 5468
rect 5409 5466 5433 5468
rect 5489 5466 5513 5468
rect 5569 5466 5575 5468
rect 5329 5414 5331 5466
rect 5511 5414 5513 5466
rect 5267 5412 5273 5414
rect 5329 5412 5353 5414
rect 5409 5412 5433 5414
rect 5489 5412 5513 5414
rect 5569 5412 5575 5414
rect 5267 5403 5575 5412
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5267 4380 5575 4389
rect 5267 4378 5273 4380
rect 5329 4378 5353 4380
rect 5409 4378 5433 4380
rect 5489 4378 5513 4380
rect 5569 4378 5575 4380
rect 5329 4326 5331 4378
rect 5511 4326 5513 4378
rect 5267 4324 5273 4326
rect 5329 4324 5353 4326
rect 5409 4324 5433 4326
rect 5489 4324 5513 4326
rect 5569 4324 5575 4326
rect 5267 4315 5575 4324
rect 5644 4078 5672 5510
rect 5736 4214 5764 5782
rect 5828 4826 5856 6938
rect 5920 6662 5948 9930
rect 6288 9722 6316 10202
rect 6656 10130 6684 10406
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6932 10010 6960 10610
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7045 10364 7353 10373
rect 7045 10362 7051 10364
rect 7107 10362 7131 10364
rect 7187 10362 7211 10364
rect 7267 10362 7291 10364
rect 7347 10362 7353 10364
rect 7107 10310 7109 10362
rect 7289 10310 7291 10362
rect 7045 10308 7051 10310
rect 7107 10308 7131 10310
rect 7187 10308 7211 10310
rect 7267 10308 7291 10310
rect 7347 10308 7353 10310
rect 7045 10299 7353 10308
rect 6460 9988 6512 9994
rect 6932 9982 7144 10010
rect 6460 9930 6512 9936
rect 6472 9722 6500 9930
rect 6828 9920 6880 9926
rect 7012 9920 7064 9926
rect 6880 9880 6960 9908
rect 6828 9862 6880 9868
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6472 8022 6500 9454
rect 6840 9382 6868 9454
rect 6932 9382 6960 9880
rect 7012 9862 7064 9868
rect 7024 9654 7052 9862
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7116 9466 7144 9982
rect 7392 9586 7420 10542
rect 7484 10062 7512 10746
rect 8128 10674 8156 13382
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8220 11150 8248 11834
rect 9483 11452 9791 11461
rect 9483 11450 9489 11452
rect 9545 11450 9569 11452
rect 9625 11450 9649 11452
rect 9705 11450 9729 11452
rect 9785 11450 9791 11452
rect 9545 11398 9547 11450
rect 9727 11398 9729 11450
rect 9483 11396 9489 11398
rect 9545 11396 9569 11398
rect 9625 11396 9649 11398
rect 9705 11396 9729 11398
rect 9785 11396 9791 11398
rect 9483 11387 9791 11396
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7668 10130 7696 10610
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 8220 10062 8248 10678
rect 8312 10538 8340 10950
rect 10143 10908 10451 10917
rect 10143 10906 10149 10908
rect 10205 10906 10229 10908
rect 10285 10906 10309 10908
rect 10365 10906 10389 10908
rect 10445 10906 10451 10908
rect 10205 10854 10207 10906
rect 10387 10854 10389 10906
rect 10143 10852 10149 10854
rect 10205 10852 10229 10854
rect 10285 10852 10309 10854
rect 10365 10852 10389 10854
rect 10445 10852 10451 10854
rect 10143 10843 10451 10852
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7705 9820 8013 9829
rect 7705 9818 7711 9820
rect 7767 9818 7791 9820
rect 7847 9818 7871 9820
rect 7927 9818 7951 9820
rect 8007 9818 8013 9820
rect 7767 9766 7769 9818
rect 7949 9766 7951 9818
rect 7705 9764 7711 9766
rect 7767 9764 7791 9766
rect 7847 9764 7871 9766
rect 7927 9764 7951 9766
rect 8007 9764 8013 9766
rect 7705 9755 8013 9764
rect 8220 9586 8248 9998
rect 8312 9926 8340 10474
rect 8588 10062 8616 10542
rect 9483 10364 9791 10373
rect 9483 10362 9489 10364
rect 9545 10362 9569 10364
rect 9625 10362 9649 10364
rect 9705 10362 9729 10364
rect 9785 10362 9791 10364
rect 9545 10310 9547 10362
rect 9727 10310 9729 10362
rect 9483 10308 9489 10310
rect 9545 10308 9569 10310
rect 9625 10308 9649 10310
rect 9705 10308 9729 10310
rect 9785 10308 9791 10310
rect 9483 10299 9791 10308
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9586 8340 9862
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8588 9518 8616 9998
rect 10143 9820 10451 9829
rect 10143 9818 10149 9820
rect 10205 9818 10229 9820
rect 10285 9818 10309 9820
rect 10365 9818 10389 9820
rect 10445 9818 10451 9820
rect 10205 9766 10207 9818
rect 10387 9766 10389 9818
rect 10143 9764 10149 9766
rect 10205 9764 10229 9766
rect 10285 9764 10309 9766
rect 10365 9764 10389 9766
rect 10445 9764 10451 9766
rect 10143 9755 10451 9764
rect 8576 9512 8628 9518
rect 7116 9438 7420 9466
rect 8576 9454 8628 9460
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6840 8090 6868 9318
rect 7045 9276 7353 9285
rect 7045 9274 7051 9276
rect 7107 9274 7131 9276
rect 7187 9274 7211 9276
rect 7267 9274 7291 9276
rect 7347 9274 7353 9276
rect 7107 9222 7109 9274
rect 7289 9222 7291 9274
rect 7045 9220 7051 9222
rect 7107 9220 7131 9222
rect 7187 9220 7211 9222
rect 7267 9220 7291 9222
rect 7347 9220 7353 9222
rect 7045 9211 7353 9220
rect 7045 8188 7353 8197
rect 7045 8186 7051 8188
rect 7107 8186 7131 8188
rect 7187 8186 7211 8188
rect 7267 8186 7291 8188
rect 7347 8186 7353 8188
rect 7107 8134 7109 8186
rect 7289 8134 7291 8186
rect 7045 8132 7051 8134
rect 7107 8132 7131 8134
rect 7187 8132 7211 8134
rect 7267 8132 7291 8134
rect 7347 8132 7353 8134
rect 7045 8123 7353 8132
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6012 6934 6040 7346
rect 6196 7342 6224 7754
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6196 6730 6224 7278
rect 6472 7274 6500 7822
rect 6564 7546 6592 7822
rect 6748 7750 6776 7958
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6748 7410 6776 7686
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6748 6798 6776 7346
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 5920 5846 5948 6598
rect 6564 5914 6592 6598
rect 6748 6390 6776 6734
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6472 5234 6500 5510
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6656 4690 6684 5714
rect 6840 5273 6868 8026
rect 7392 8004 7420 9438
rect 8588 9178 8616 9454
rect 9483 9276 9791 9285
rect 9483 9274 9489 9276
rect 9545 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9791 9276
rect 9545 9222 9547 9274
rect 9727 9222 9729 9274
rect 9483 9220 9489 9222
rect 9545 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9791 9222
rect 9483 9211 9791 9220
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9128 8968 9180 8974
rect 10508 8968 10560 8974
rect 9128 8910 9180 8916
rect 10506 8936 10508 8945
rect 10560 8936 10562 8945
rect 7705 8732 8013 8741
rect 7705 8730 7711 8732
rect 7767 8730 7791 8732
rect 7847 8730 7871 8732
rect 7927 8730 7951 8732
rect 8007 8730 8013 8732
rect 7767 8678 7769 8730
rect 7949 8678 7951 8730
rect 7705 8676 7711 8678
rect 7767 8676 7791 8678
rect 7847 8676 7871 8678
rect 7927 8676 7951 8678
rect 8007 8676 8013 8678
rect 7705 8667 8013 8676
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 7300 7976 7420 8004
rect 8024 8016 8076 8022
rect 7104 7880 7156 7886
rect 7024 7840 7104 7868
rect 7024 7342 7052 7840
rect 7300 7868 7328 7976
rect 8076 7964 8248 7970
rect 8024 7958 8248 7964
rect 8036 7954 8248 7958
rect 8036 7948 8260 7954
rect 8036 7942 8208 7948
rect 8208 7890 8260 7896
rect 8588 7886 8616 8298
rect 7156 7840 7328 7868
rect 7380 7880 7432 7886
rect 7104 7822 7156 7828
rect 7380 7822 7432 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7410 7144 7686
rect 7392 7546 7420 7822
rect 7705 7644 8013 7653
rect 7705 7642 7711 7644
rect 7767 7642 7791 7644
rect 7847 7642 7871 7644
rect 7927 7642 7951 7644
rect 8007 7642 8013 7644
rect 7767 7590 7769 7642
rect 7949 7590 7951 7642
rect 7705 7588 7711 7590
rect 7767 7588 7791 7590
rect 7847 7588 7871 7590
rect 7927 7588 7951 7590
rect 8007 7588 8013 7590
rect 7705 7579 8013 7588
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 8404 7410 8432 7822
rect 8680 7818 8708 8434
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8680 7546 8708 7754
rect 8864 7750 8892 7890
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8864 7478 8892 7686
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7045 7100 7353 7109
rect 7045 7098 7051 7100
rect 7107 7098 7131 7100
rect 7187 7098 7211 7100
rect 7267 7098 7291 7100
rect 7347 7098 7353 7100
rect 7107 7046 7109 7098
rect 7289 7046 7291 7098
rect 7045 7044 7051 7046
rect 7107 7044 7131 7046
rect 7187 7044 7211 7046
rect 7267 7044 7291 7046
rect 7347 7044 7353 7046
rect 7045 7035 7353 7044
rect 8588 7002 8616 7346
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8864 6866 8892 7414
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7045 6012 7353 6021
rect 7045 6010 7051 6012
rect 7107 6010 7131 6012
rect 7187 6010 7211 6012
rect 7267 6010 7291 6012
rect 7347 6010 7353 6012
rect 7107 5958 7109 6010
rect 7289 5958 7291 6010
rect 7045 5956 7051 5958
rect 7107 5956 7131 5958
rect 7187 5956 7211 5958
rect 7267 5956 7291 5958
rect 7347 5956 7353 5958
rect 7045 5947 7353 5956
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6932 5710 6960 5782
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 6826 5264 6882 5273
rect 6826 5199 6882 5208
rect 6736 5160 6788 5166
rect 6932 5114 6960 5646
rect 7208 5370 7236 5646
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6736 5102 6788 5108
rect 6748 4826 6776 5102
rect 6840 5086 6960 5114
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 4172 3998 4384 4026
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 4436 4004 4488 4010
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 3514 3632 3570 3641
rect 4172 3602 4200 3998
rect 4436 3946 4488 3952
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 3514 3567 3516 3576
rect 3568 3567 3570 3576
rect 4160 3596 4212 3602
rect 3516 3538 3568 3544
rect 4160 3538 4212 3544
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 2056 3194 2084 3470
rect 2228 3392 2280 3398
rect 2792 3380 2820 3470
rect 2228 3334 2280 3340
rect 2700 3352 2820 3380
rect 3240 3392 3292 3398
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2240 3058 2268 3334
rect 2700 3176 2728 3352
rect 3240 3334 3292 3340
rect 2829 3292 3137 3301
rect 2829 3290 2835 3292
rect 2891 3290 2915 3292
rect 2971 3290 2995 3292
rect 3051 3290 3075 3292
rect 3131 3290 3137 3292
rect 2891 3238 2893 3290
rect 3073 3238 3075 3290
rect 2829 3236 2835 3238
rect 2891 3236 2915 3238
rect 2971 3236 2995 3238
rect 3051 3236 3075 3238
rect 3131 3236 3137 3238
rect 2829 3227 3137 3236
rect 2780 3188 2832 3194
rect 2700 3148 2780 3176
rect 2780 3130 2832 3136
rect 3252 3126 3280 3334
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 3344 2922 3372 3470
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3436 3194 3464 3402
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4066 3088 4122 3097
rect 4066 3023 4068 3032
rect 4120 3023 4122 3032
rect 4068 2994 4120 3000
rect 4172 2990 4200 3538
rect 4356 3126 4384 3878
rect 4448 3398 4476 3946
rect 5644 3942 5672 4014
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 4540 3670 4568 3878
rect 4607 3836 4915 3845
rect 4607 3834 4613 3836
rect 4669 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4915 3836
rect 4669 3782 4671 3834
rect 4851 3782 4853 3834
rect 4607 3780 4613 3782
rect 4669 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4915 3782
rect 4607 3771 4915 3780
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4632 3602 4660 3674
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 5000 3534 5028 3878
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 2169 2748 2477 2757
rect 2169 2746 2175 2748
rect 2231 2746 2255 2748
rect 2311 2746 2335 2748
rect 2391 2746 2415 2748
rect 2471 2746 2477 2748
rect 2231 2694 2233 2746
rect 2413 2694 2415 2746
rect 2169 2692 2175 2694
rect 2231 2692 2255 2694
rect 2311 2692 2335 2694
rect 2391 2692 2415 2694
rect 2471 2692 2477 2694
rect 2169 2683 2477 2692
rect 4172 2650 4200 2926
rect 4356 2922 4384 3062
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4448 2650 4476 3334
rect 4540 3194 4568 3470
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 5000 3058 5028 3470
rect 5092 3194 5120 3470
rect 5184 3194 5212 3538
rect 5267 3292 5575 3301
rect 5267 3290 5273 3292
rect 5329 3290 5353 3292
rect 5409 3290 5433 3292
rect 5489 3290 5513 3292
rect 5569 3290 5575 3292
rect 5329 3238 5331 3290
rect 5511 3238 5513 3290
rect 5267 3236 5273 3238
rect 5329 3236 5353 3238
rect 5409 3236 5433 3238
rect 5489 3236 5513 3238
rect 5569 3236 5575 3238
rect 5267 3227 5575 3236
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5644 2854 5672 3878
rect 5736 3534 5764 4150
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 4607 2748 4915 2757
rect 4607 2746 4613 2748
rect 4669 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4915 2748
rect 4669 2694 4671 2746
rect 4851 2694 4853 2746
rect 4607 2692 4613 2694
rect 4669 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4915 2694
rect 4607 2683 4915 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5736 2446 5764 3334
rect 5828 3126 5856 3878
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6472 2650 6500 4558
rect 6656 3738 6684 4626
rect 6748 4214 6776 4762
rect 6840 4622 6868 5086
rect 7300 5030 7328 5850
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6656 3466 6684 3674
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6932 2446 6960 4966
rect 7045 4924 7353 4933
rect 7045 4922 7051 4924
rect 7107 4922 7131 4924
rect 7187 4922 7211 4924
rect 7267 4922 7291 4924
rect 7347 4922 7353 4924
rect 7107 4870 7109 4922
rect 7289 4870 7291 4922
rect 7045 4868 7051 4870
rect 7107 4868 7131 4870
rect 7187 4868 7211 4870
rect 7267 4868 7291 4870
rect 7347 4868 7353 4870
rect 7045 4859 7353 4868
rect 7392 4690 7420 6666
rect 7705 6556 8013 6565
rect 7705 6554 7711 6556
rect 7767 6554 7791 6556
rect 7847 6554 7871 6556
rect 7927 6554 7951 6556
rect 8007 6554 8013 6556
rect 7767 6502 7769 6554
rect 7949 6502 7951 6554
rect 7705 6500 7711 6502
rect 7767 6500 7791 6502
rect 7847 6500 7871 6502
rect 7927 6500 7951 6502
rect 8007 6500 8013 6502
rect 7705 6491 8013 6500
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7668 5710 7696 5850
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 8024 5636 8076 5642
rect 8076 5596 8156 5624
rect 8024 5578 8076 5584
rect 7484 5370 7512 5578
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7470 5264 7526 5273
rect 7470 5199 7472 5208
rect 7524 5199 7526 5208
rect 7472 5170 7524 5176
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 4214 7420 4626
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7045 3836 7353 3845
rect 7045 3834 7051 3836
rect 7107 3834 7131 3836
rect 7187 3834 7211 3836
rect 7267 3834 7291 3836
rect 7347 3834 7353 3836
rect 7107 3782 7109 3834
rect 7289 3782 7291 3834
rect 7045 3780 7051 3782
rect 7107 3780 7131 3782
rect 7187 3780 7211 3782
rect 7267 3780 7291 3782
rect 7347 3780 7353 3782
rect 7045 3771 7353 3780
rect 7484 3641 7512 5170
rect 7576 4826 7604 5510
rect 7705 5468 8013 5477
rect 7705 5466 7711 5468
rect 7767 5466 7791 5468
rect 7847 5466 7871 5468
rect 7927 5466 7951 5468
rect 8007 5466 8013 5468
rect 7767 5414 7769 5466
rect 7949 5414 7951 5466
rect 7705 5412 7711 5414
rect 7767 5412 7791 5414
rect 7847 5412 7871 5414
rect 7927 5412 7951 5414
rect 8007 5412 8013 5414
rect 7705 5403 8013 5412
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 5030 7696 5170
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7668 4706 7696 4966
rect 7576 4678 7696 4706
rect 7470 3632 7526 3641
rect 7380 3596 7432 3602
rect 7470 3567 7526 3576
rect 7380 3538 7432 3544
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7024 3194 7052 3334
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7116 3097 7144 3334
rect 7392 3194 7420 3538
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7484 3126 7512 3567
rect 7576 3534 7604 4678
rect 8024 4616 8076 4622
rect 8128 4604 8156 5596
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 5302 8248 5510
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8076 4576 8156 4604
rect 8024 4558 8076 4564
rect 8220 4486 8248 5238
rect 8404 5234 8432 6190
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8588 5642 8616 5850
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8588 5234 8616 5578
rect 8772 5574 8800 6258
rect 8956 5914 8984 8910
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8498 9076 8774
rect 9140 8634 9168 8910
rect 9404 8900 9456 8906
rect 10506 8871 10562 8880
rect 9404 8842 9456 8848
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9312 8424 9364 8430
rect 9232 8384 9312 8412
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8022 9076 8230
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9048 7562 9076 7958
rect 9232 7818 9260 8384
rect 9312 8366 9364 8372
rect 9416 8090 9444 8842
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9876 8498 9904 8774
rect 9968 8566 9996 8774
rect 10143 8732 10451 8741
rect 10143 8730 10149 8732
rect 10205 8730 10229 8732
rect 10285 8730 10309 8732
rect 10365 8730 10389 8732
rect 10445 8730 10451 8732
rect 10205 8678 10207 8730
rect 10387 8678 10389 8730
rect 10143 8676 10149 8678
rect 10205 8676 10229 8678
rect 10285 8676 10309 8678
rect 10365 8676 10389 8678
rect 10445 8676 10451 8678
rect 10143 8667 10451 8676
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 8294 9536 8366
rect 9600 8294 9628 8434
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9483 8188 9791 8197
rect 9483 8186 9489 8188
rect 9545 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9791 8188
rect 9545 8134 9547 8186
rect 9727 8134 9729 8186
rect 9483 8132 9489 8134
rect 9545 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9791 8134
rect 9483 8123 9791 8132
rect 9876 8090 9904 8434
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9496 7880 9548 7886
rect 9416 7828 9496 7834
rect 9416 7822 9548 7828
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9312 7812 9364 7818
rect 9416 7806 9536 7822
rect 9416 7800 9444 7806
rect 9364 7772 9444 7800
rect 9312 7754 9364 7760
rect 9048 7534 9168 7562
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 6780 9076 7346
rect 9140 7274 9168 7534
rect 9232 7410 9260 7754
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7546 9536 7686
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9876 7478 9904 8026
rect 9968 7886 9996 8230
rect 10244 8022 10272 8434
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10506 8256 10562 8265
rect 10506 8191 10562 8200
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10520 7886 10548 8191
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9483 7100 9791 7109
rect 9483 7098 9489 7100
rect 9545 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9791 7100
rect 9545 7046 9547 7098
rect 9727 7046 9729 7098
rect 9483 7044 9489 7046
rect 9545 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9791 7046
rect 9483 7035 9791 7044
rect 9876 6934 9904 7278
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9968 6798 9996 7822
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 6866 10088 7754
rect 10143 7644 10451 7653
rect 10143 7642 10149 7644
rect 10205 7642 10229 7644
rect 10285 7642 10309 7644
rect 10365 7642 10389 7644
rect 10445 7642 10451 7644
rect 10205 7590 10207 7642
rect 10387 7590 10389 7642
rect 10143 7588 10149 7590
rect 10205 7588 10229 7590
rect 10285 7588 10309 7590
rect 10365 7588 10389 7590
rect 10445 7588 10451 7590
rect 10143 7579 10451 7588
rect 10704 7585 10732 8298
rect 10690 7576 10746 7585
rect 10690 7511 10746 7520
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10244 6798 10272 7346
rect 10428 6905 10456 7346
rect 10414 6896 10470 6905
rect 10414 6831 10470 6840
rect 9128 6792 9180 6798
rect 9048 6752 9128 6780
rect 9128 6734 9180 6740
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9140 6458 9168 6734
rect 9232 6662 9260 6734
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8404 4706 8432 5170
rect 8772 5098 8800 5510
rect 8864 5098 8892 5646
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8312 4690 8432 4706
rect 8956 4690 8984 5646
rect 8300 4684 8432 4690
rect 8352 4678 8432 4684
rect 8300 4626 8352 4632
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7705 4380 8013 4389
rect 7705 4378 7711 4380
rect 7767 4378 7791 4380
rect 7847 4378 7871 4380
rect 7927 4378 7951 4380
rect 8007 4378 8013 4380
rect 7767 4326 7769 4378
rect 7949 4326 7951 4378
rect 7705 4324 7711 4326
rect 7767 4324 7791 4326
rect 7847 4324 7871 4326
rect 7927 4324 7951 4326
rect 8007 4324 8013 4326
rect 7705 4315 8013 4324
rect 8312 3534 8340 4490
rect 8404 3670 8432 4678
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 4146 8984 4626
rect 9048 4622 9076 6258
rect 9324 5234 9352 6258
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9416 5710 9444 6122
rect 9483 6012 9791 6021
rect 9483 6010 9489 6012
rect 9545 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9791 6012
rect 9545 5958 9547 6010
rect 9727 5958 9729 6010
rect 9483 5956 9489 5958
rect 9545 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9791 5958
rect 9483 5947 9791 5956
rect 9968 5846 9996 6734
rect 10143 6556 10451 6565
rect 10143 6554 10149 6556
rect 10205 6554 10229 6556
rect 10285 6554 10309 6556
rect 10365 6554 10389 6556
rect 10445 6554 10451 6556
rect 10205 6502 10207 6554
rect 10387 6502 10389 6554
rect 10143 6500 10149 6502
rect 10205 6500 10229 6502
rect 10285 6500 10309 6502
rect 10365 6500 10389 6502
rect 10445 6500 10451 6502
rect 10143 6491 10451 6500
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10048 6248 10100 6254
rect 10428 6225 10456 6258
rect 10048 6190 10100 6196
rect 10414 6216 10470 6225
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 4690 9352 5034
rect 9483 4924 9791 4933
rect 9483 4922 9489 4924
rect 9545 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9791 4924
rect 9545 4870 9547 4922
rect 9727 4870 9729 4922
rect 9483 4868 9489 4870
rect 9545 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9791 4870
rect 9483 4859 9791 4868
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8864 3602 8892 4014
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 9140 3534 9168 3674
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7472 3120 7524 3126
rect 7102 3088 7158 3097
rect 7472 3062 7524 3068
rect 7576 3058 7604 3334
rect 7705 3292 8013 3301
rect 7705 3290 7711 3292
rect 7767 3290 7791 3292
rect 7847 3290 7871 3292
rect 7927 3290 7951 3292
rect 8007 3290 8013 3292
rect 7767 3238 7769 3290
rect 7949 3238 7951 3290
rect 7705 3236 7711 3238
rect 7767 3236 7791 3238
rect 7847 3236 7871 3238
rect 7927 3236 7951 3238
rect 8007 3236 8013 3238
rect 7705 3227 8013 3236
rect 7102 3023 7158 3032
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 8404 2990 8432 3470
rect 8496 3058 8524 3470
rect 8956 3398 8984 3470
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3194 8984 3334
rect 9324 3194 9352 3470
rect 9416 3466 9444 3878
rect 9483 3836 9791 3845
rect 9483 3834 9489 3836
rect 9545 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9791 3836
rect 9545 3782 9547 3834
rect 9727 3782 9729 3834
rect 9483 3780 9489 3782
rect 9545 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9791 3782
rect 9483 3771 9791 3780
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9404 3460 9456 3466
rect 9404 3402 9456 3408
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8496 2854 8524 2994
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 7045 2748 7353 2757
rect 7045 2746 7051 2748
rect 7107 2746 7131 2748
rect 7187 2746 7211 2748
rect 7267 2746 7291 2748
rect 7347 2746 7353 2748
rect 7107 2694 7109 2746
rect 7289 2694 7291 2746
rect 7045 2692 7051 2694
rect 7107 2692 7131 2694
rect 7187 2692 7211 2694
rect 7267 2692 7291 2694
rect 7347 2692 7353 2694
rect 7045 2683 7353 2692
rect 7852 2446 7880 2790
rect 8680 2650 8708 3062
rect 9416 3058 9444 3402
rect 9692 3194 9720 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9600 3074 9628 3130
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9508 2990 9536 3062
rect 9600 3058 9812 3074
rect 9876 3058 9904 4082
rect 9968 3126 9996 4082
rect 10060 3738 10088 6190
rect 10414 6151 10470 6160
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10612 5545 10640 5646
rect 10598 5536 10654 5545
rect 10143 5468 10451 5477
rect 10598 5471 10654 5480
rect 10143 5466 10149 5468
rect 10205 5466 10229 5468
rect 10285 5466 10309 5468
rect 10365 5466 10389 5468
rect 10445 5466 10451 5468
rect 10205 5414 10207 5466
rect 10387 5414 10389 5466
rect 10143 5412 10149 5414
rect 10205 5412 10229 5414
rect 10285 5412 10309 5414
rect 10365 5412 10389 5414
rect 10445 5412 10451 5414
rect 10143 5403 10451 5412
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10520 4865 10548 5170
rect 10506 4856 10562 4865
rect 10506 4791 10562 4800
rect 10143 4380 10451 4389
rect 10143 4378 10149 4380
rect 10205 4378 10229 4380
rect 10285 4378 10309 4380
rect 10365 4378 10389 4380
rect 10445 4378 10451 4380
rect 10205 4326 10207 4378
rect 10387 4326 10389 4378
rect 10143 4324 10149 4326
rect 10205 4324 10229 4326
rect 10285 4324 10309 4326
rect 10365 4324 10389 4326
rect 10445 4324 10451 4326
rect 10143 4315 10451 4324
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10143 3292 10451 3301
rect 10143 3290 10149 3292
rect 10205 3290 10229 3292
rect 10285 3290 10309 3292
rect 10365 3290 10389 3292
rect 10445 3290 10451 3292
rect 10205 3238 10207 3290
rect 10387 3238 10389 3290
rect 10143 3236 10149 3238
rect 10205 3236 10229 3238
rect 10285 3236 10309 3238
rect 10365 3236 10389 3238
rect 10445 3236 10451 3238
rect 10143 3227 10451 3236
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9600 3052 9824 3058
rect 9600 3046 9772 3052
rect 9772 2994 9824 3000
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9496 2984 9548 2990
rect 9416 2932 9496 2938
rect 9416 2926 9548 2932
rect 9784 2938 9812 2994
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9416 2910 9536 2926
rect 9784 2910 9904 2938
rect 9232 2650 9260 2858
rect 9416 2774 9444 2910
rect 9324 2746 9444 2774
rect 9483 2748 9791 2757
rect 9483 2746 9489 2748
rect 9545 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9791 2748
rect 9324 2650 9352 2746
rect 9545 2694 9547 2746
rect 9727 2694 9729 2746
rect 9483 2692 9489 2694
rect 9545 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9791 2694
rect 9483 2683 9791 2692
rect 9876 2650 9904 2910
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 2829 2204 3137 2213
rect 2829 2202 2835 2204
rect 2891 2202 2915 2204
rect 2971 2202 2995 2204
rect 3051 2202 3075 2204
rect 3131 2202 3137 2204
rect 2891 2150 2893 2202
rect 3073 2150 3075 2202
rect 2829 2148 2835 2150
rect 2891 2148 2915 2150
rect 2971 2148 2995 2150
rect 3051 2148 3075 2150
rect 3131 2148 3137 2150
rect 2829 2139 3137 2148
rect 3896 800 3924 2382
rect 4540 800 4568 2382
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 5184 800 5212 2314
rect 5267 2204 5575 2213
rect 5267 2202 5273 2204
rect 5329 2202 5353 2204
rect 5409 2202 5433 2204
rect 5489 2202 5513 2204
rect 5569 2202 5575 2204
rect 5329 2150 5331 2202
rect 5511 2150 5513 2202
rect 5267 2148 5273 2150
rect 5329 2148 5353 2150
rect 5409 2148 5433 2150
rect 5489 2148 5513 2150
rect 5569 2148 5575 2150
rect 5267 2139 5575 2148
rect 6472 800 6500 2382
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7116 800 7144 2246
rect 7576 1170 7604 2246
rect 7705 2204 8013 2213
rect 7705 2202 7711 2204
rect 7767 2202 7791 2204
rect 7847 2202 7871 2204
rect 7927 2202 7951 2204
rect 8007 2202 8013 2204
rect 7767 2150 7769 2202
rect 7949 2150 7951 2202
rect 7705 2148 7711 2150
rect 7767 2148 7791 2150
rect 7847 2148 7871 2150
rect 7927 2148 7951 2150
rect 8007 2148 8013 2150
rect 7705 2139 8013 2148
rect 7576 1142 7788 1170
rect 7760 800 7788 1142
rect 8404 800 8432 2382
rect 9048 800 9076 2382
rect 9692 800 9720 2382
rect 10143 2204 10451 2213
rect 10143 2202 10149 2204
rect 10205 2202 10229 2204
rect 10285 2202 10309 2204
rect 10365 2202 10389 2204
rect 10445 2202 10451 2204
rect 10205 2150 10207 2202
rect 10387 2150 10389 2202
rect 10143 2148 10149 2150
rect 10205 2148 10229 2150
rect 10285 2148 10309 2150
rect 10365 2148 10389 2150
rect 10445 2148 10451 2150
rect 10143 2139 10451 2148
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
<< via2 >>
rect 2175 11450 2231 11452
rect 2255 11450 2311 11452
rect 2335 11450 2391 11452
rect 2415 11450 2471 11452
rect 2175 11398 2221 11450
rect 2221 11398 2231 11450
rect 2255 11398 2285 11450
rect 2285 11398 2297 11450
rect 2297 11398 2311 11450
rect 2335 11398 2349 11450
rect 2349 11398 2361 11450
rect 2361 11398 2391 11450
rect 2415 11398 2425 11450
rect 2425 11398 2471 11450
rect 2175 11396 2231 11398
rect 2255 11396 2311 11398
rect 2335 11396 2391 11398
rect 2415 11396 2471 11398
rect 4613 11450 4669 11452
rect 4693 11450 4749 11452
rect 4773 11450 4829 11452
rect 4853 11450 4909 11452
rect 4613 11398 4659 11450
rect 4659 11398 4669 11450
rect 4693 11398 4723 11450
rect 4723 11398 4735 11450
rect 4735 11398 4749 11450
rect 4773 11398 4787 11450
rect 4787 11398 4799 11450
rect 4799 11398 4829 11450
rect 4853 11398 4863 11450
rect 4863 11398 4909 11450
rect 4613 11396 4669 11398
rect 4693 11396 4749 11398
rect 4773 11396 4829 11398
rect 4853 11396 4909 11398
rect 7051 11450 7107 11452
rect 7131 11450 7187 11452
rect 7211 11450 7267 11452
rect 7291 11450 7347 11452
rect 7051 11398 7097 11450
rect 7097 11398 7107 11450
rect 7131 11398 7161 11450
rect 7161 11398 7173 11450
rect 7173 11398 7187 11450
rect 7211 11398 7225 11450
rect 7225 11398 7237 11450
rect 7237 11398 7267 11450
rect 7291 11398 7301 11450
rect 7301 11398 7347 11450
rect 7051 11396 7107 11398
rect 7131 11396 7187 11398
rect 7211 11396 7267 11398
rect 7291 11396 7347 11398
rect 2835 10906 2891 10908
rect 2915 10906 2971 10908
rect 2995 10906 3051 10908
rect 3075 10906 3131 10908
rect 2835 10854 2881 10906
rect 2881 10854 2891 10906
rect 2915 10854 2945 10906
rect 2945 10854 2957 10906
rect 2957 10854 2971 10906
rect 2995 10854 3009 10906
rect 3009 10854 3021 10906
rect 3021 10854 3051 10906
rect 3075 10854 3085 10906
rect 3085 10854 3131 10906
rect 2835 10852 2891 10854
rect 2915 10852 2971 10854
rect 2995 10852 3051 10854
rect 3075 10852 3131 10854
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 846 9016 902 9072
rect 2175 10362 2231 10364
rect 2255 10362 2311 10364
rect 2335 10362 2391 10364
rect 2415 10362 2471 10364
rect 2175 10310 2221 10362
rect 2221 10310 2231 10362
rect 2255 10310 2285 10362
rect 2285 10310 2297 10362
rect 2297 10310 2311 10362
rect 2335 10310 2349 10362
rect 2349 10310 2361 10362
rect 2361 10310 2391 10362
rect 2415 10310 2425 10362
rect 2425 10310 2471 10362
rect 2175 10308 2231 10310
rect 2255 10308 2311 10310
rect 2335 10308 2391 10310
rect 2415 10308 2471 10310
rect 1490 8200 1546 8256
rect 846 7404 902 7440
rect 2835 9818 2891 9820
rect 2915 9818 2971 9820
rect 2995 9818 3051 9820
rect 3075 9818 3131 9820
rect 2835 9766 2881 9818
rect 2881 9766 2891 9818
rect 2915 9766 2945 9818
rect 2945 9766 2957 9818
rect 2957 9766 2971 9818
rect 2995 9766 3009 9818
rect 3009 9766 3021 9818
rect 3021 9766 3051 9818
rect 3075 9766 3085 9818
rect 3085 9766 3131 9818
rect 2835 9764 2891 9766
rect 2915 9764 2971 9766
rect 2995 9764 3051 9766
rect 3075 9764 3131 9766
rect 5273 10906 5329 10908
rect 5353 10906 5409 10908
rect 5433 10906 5489 10908
rect 5513 10906 5569 10908
rect 5273 10854 5319 10906
rect 5319 10854 5329 10906
rect 5353 10854 5383 10906
rect 5383 10854 5395 10906
rect 5395 10854 5409 10906
rect 5433 10854 5447 10906
rect 5447 10854 5459 10906
rect 5459 10854 5489 10906
rect 5513 10854 5523 10906
rect 5523 10854 5569 10906
rect 5273 10852 5329 10854
rect 5353 10852 5409 10854
rect 5433 10852 5489 10854
rect 5513 10852 5569 10854
rect 7711 10906 7767 10908
rect 7791 10906 7847 10908
rect 7871 10906 7927 10908
rect 7951 10906 8007 10908
rect 7711 10854 7757 10906
rect 7757 10854 7767 10906
rect 7791 10854 7821 10906
rect 7821 10854 7833 10906
rect 7833 10854 7847 10906
rect 7871 10854 7885 10906
rect 7885 10854 7897 10906
rect 7897 10854 7927 10906
rect 7951 10854 7961 10906
rect 7961 10854 8007 10906
rect 7711 10852 7767 10854
rect 7791 10852 7847 10854
rect 7871 10852 7927 10854
rect 7951 10852 8007 10854
rect 4613 10362 4669 10364
rect 4693 10362 4749 10364
rect 4773 10362 4829 10364
rect 4853 10362 4909 10364
rect 4613 10310 4659 10362
rect 4659 10310 4669 10362
rect 4693 10310 4723 10362
rect 4723 10310 4735 10362
rect 4735 10310 4749 10362
rect 4773 10310 4787 10362
rect 4787 10310 4799 10362
rect 4799 10310 4829 10362
rect 4853 10310 4863 10362
rect 4863 10310 4909 10362
rect 4613 10308 4669 10310
rect 4693 10308 4749 10310
rect 4773 10308 4829 10310
rect 4853 10308 4909 10310
rect 2175 9274 2231 9276
rect 2255 9274 2311 9276
rect 2335 9274 2391 9276
rect 2415 9274 2471 9276
rect 2175 9222 2221 9274
rect 2221 9222 2231 9274
rect 2255 9222 2285 9274
rect 2285 9222 2297 9274
rect 2297 9222 2311 9274
rect 2335 9222 2349 9274
rect 2349 9222 2361 9274
rect 2361 9222 2391 9274
rect 2415 9222 2425 9274
rect 2425 9222 2471 9274
rect 2175 9220 2231 9222
rect 2255 9220 2311 9222
rect 2335 9220 2391 9222
rect 2415 9220 2471 9222
rect 2835 8730 2891 8732
rect 2915 8730 2971 8732
rect 2995 8730 3051 8732
rect 3075 8730 3131 8732
rect 2835 8678 2881 8730
rect 2881 8678 2891 8730
rect 2915 8678 2945 8730
rect 2945 8678 2957 8730
rect 2957 8678 2971 8730
rect 2995 8678 3009 8730
rect 3009 8678 3021 8730
rect 3021 8678 3051 8730
rect 3075 8678 3085 8730
rect 3085 8678 3131 8730
rect 2835 8676 2891 8678
rect 2915 8676 2971 8678
rect 2995 8676 3051 8678
rect 3075 8676 3131 8678
rect 846 7384 848 7404
rect 848 7384 900 7404
rect 900 7384 902 7404
rect 2175 8186 2231 8188
rect 2255 8186 2311 8188
rect 2335 8186 2391 8188
rect 2415 8186 2471 8188
rect 2175 8134 2221 8186
rect 2221 8134 2231 8186
rect 2255 8134 2285 8186
rect 2285 8134 2297 8186
rect 2297 8134 2311 8186
rect 2335 8134 2349 8186
rect 2349 8134 2361 8186
rect 2361 8134 2391 8186
rect 2415 8134 2425 8186
rect 2425 8134 2471 8186
rect 2175 8132 2231 8134
rect 2255 8132 2311 8134
rect 2335 8132 2391 8134
rect 2415 8132 2471 8134
rect 5273 9818 5329 9820
rect 5353 9818 5409 9820
rect 5433 9818 5489 9820
rect 5513 9818 5569 9820
rect 5273 9766 5319 9818
rect 5319 9766 5329 9818
rect 5353 9766 5383 9818
rect 5383 9766 5395 9818
rect 5395 9766 5409 9818
rect 5433 9766 5447 9818
rect 5447 9766 5459 9818
rect 5459 9766 5489 9818
rect 5513 9766 5523 9818
rect 5523 9766 5569 9818
rect 5273 9764 5329 9766
rect 5353 9764 5409 9766
rect 5433 9764 5489 9766
rect 5513 9764 5569 9766
rect 4613 9274 4669 9276
rect 4693 9274 4749 9276
rect 4773 9274 4829 9276
rect 4853 9274 4909 9276
rect 4613 9222 4659 9274
rect 4659 9222 4669 9274
rect 4693 9222 4723 9274
rect 4723 9222 4735 9274
rect 4735 9222 4749 9274
rect 4773 9222 4787 9274
rect 4787 9222 4799 9274
rect 4799 9222 4829 9274
rect 4853 9222 4863 9274
rect 4863 9222 4909 9274
rect 4613 9220 4669 9222
rect 4693 9220 4749 9222
rect 4773 9220 4829 9222
rect 4853 9220 4909 9222
rect 2835 7642 2891 7644
rect 2915 7642 2971 7644
rect 2995 7642 3051 7644
rect 3075 7642 3131 7644
rect 2835 7590 2881 7642
rect 2881 7590 2891 7642
rect 2915 7590 2945 7642
rect 2945 7590 2957 7642
rect 2957 7590 2971 7642
rect 2995 7590 3009 7642
rect 3009 7590 3021 7642
rect 3021 7590 3051 7642
rect 3075 7590 3085 7642
rect 3085 7590 3131 7642
rect 2835 7588 2891 7590
rect 2915 7588 2971 7590
rect 2995 7588 3051 7590
rect 3075 7588 3131 7590
rect 2175 7098 2231 7100
rect 2255 7098 2311 7100
rect 2335 7098 2391 7100
rect 2415 7098 2471 7100
rect 2175 7046 2221 7098
rect 2221 7046 2231 7098
rect 2255 7046 2285 7098
rect 2285 7046 2297 7098
rect 2297 7046 2311 7098
rect 2335 7046 2349 7098
rect 2349 7046 2361 7098
rect 2361 7046 2391 7098
rect 2415 7046 2425 7098
rect 2425 7046 2471 7098
rect 2175 7044 2231 7046
rect 2255 7044 2311 7046
rect 2335 7044 2391 7046
rect 2415 7044 2471 7046
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 2835 6554 2891 6556
rect 2915 6554 2971 6556
rect 2995 6554 3051 6556
rect 3075 6554 3131 6556
rect 2835 6502 2881 6554
rect 2881 6502 2891 6554
rect 2915 6502 2945 6554
rect 2945 6502 2957 6554
rect 2957 6502 2971 6554
rect 2995 6502 3009 6554
rect 3009 6502 3021 6554
rect 3021 6502 3051 6554
rect 3075 6502 3085 6554
rect 3085 6502 3131 6554
rect 2835 6500 2891 6502
rect 2915 6500 2971 6502
rect 2995 6500 3051 6502
rect 3075 6500 3131 6502
rect 2175 6010 2231 6012
rect 2255 6010 2311 6012
rect 2335 6010 2391 6012
rect 2415 6010 2471 6012
rect 2175 5958 2221 6010
rect 2221 5958 2231 6010
rect 2255 5958 2285 6010
rect 2285 5958 2297 6010
rect 2297 5958 2311 6010
rect 2335 5958 2349 6010
rect 2349 5958 2361 6010
rect 2361 5958 2391 6010
rect 2415 5958 2425 6010
rect 2425 5958 2471 6010
rect 2175 5956 2231 5958
rect 2255 5956 2311 5958
rect 2335 5956 2391 5958
rect 2415 5956 2471 5958
rect 1306 5480 1362 5536
rect 846 4664 902 4720
rect 846 3596 902 3632
rect 2175 4922 2231 4924
rect 2255 4922 2311 4924
rect 2335 4922 2391 4924
rect 2415 4922 2471 4924
rect 2175 4870 2221 4922
rect 2221 4870 2231 4922
rect 2255 4870 2285 4922
rect 2285 4870 2297 4922
rect 2297 4870 2311 4922
rect 2335 4870 2349 4922
rect 2349 4870 2361 4922
rect 2361 4870 2391 4922
rect 2415 4870 2425 4922
rect 2425 4870 2471 4922
rect 2175 4868 2231 4870
rect 2255 4868 2311 4870
rect 2335 4868 2391 4870
rect 2415 4868 2471 4870
rect 2175 3834 2231 3836
rect 2255 3834 2311 3836
rect 2335 3834 2391 3836
rect 2415 3834 2471 3836
rect 2175 3782 2221 3834
rect 2221 3782 2231 3834
rect 2255 3782 2285 3834
rect 2285 3782 2297 3834
rect 2297 3782 2311 3834
rect 2335 3782 2349 3834
rect 2349 3782 2361 3834
rect 2361 3782 2391 3834
rect 2415 3782 2425 3834
rect 2425 3782 2471 3834
rect 2175 3780 2231 3782
rect 2255 3780 2311 3782
rect 2335 3780 2391 3782
rect 2415 3780 2471 3782
rect 2835 5466 2891 5468
rect 2915 5466 2971 5468
rect 2995 5466 3051 5468
rect 3075 5466 3131 5468
rect 2835 5414 2881 5466
rect 2881 5414 2891 5466
rect 2915 5414 2945 5466
rect 2945 5414 2957 5466
rect 2957 5414 2971 5466
rect 2995 5414 3009 5466
rect 3009 5414 3021 5466
rect 3021 5414 3051 5466
rect 3075 5414 3085 5466
rect 3085 5414 3131 5466
rect 2835 5412 2891 5414
rect 2915 5412 2971 5414
rect 2995 5412 3051 5414
rect 3075 5412 3131 5414
rect 4613 8186 4669 8188
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4613 8134 4659 8186
rect 4659 8134 4669 8186
rect 4693 8134 4723 8186
rect 4723 8134 4735 8186
rect 4735 8134 4749 8186
rect 4773 8134 4787 8186
rect 4787 8134 4799 8186
rect 4799 8134 4829 8186
rect 4853 8134 4863 8186
rect 4863 8134 4909 8186
rect 4613 8132 4669 8134
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 5273 8730 5329 8732
rect 5353 8730 5409 8732
rect 5433 8730 5489 8732
rect 5513 8730 5569 8732
rect 5273 8678 5319 8730
rect 5319 8678 5329 8730
rect 5353 8678 5383 8730
rect 5383 8678 5395 8730
rect 5395 8678 5409 8730
rect 5433 8678 5447 8730
rect 5447 8678 5459 8730
rect 5459 8678 5489 8730
rect 5513 8678 5523 8730
rect 5523 8678 5569 8730
rect 5273 8676 5329 8678
rect 5353 8676 5409 8678
rect 5433 8676 5489 8678
rect 5513 8676 5569 8678
rect 5273 7642 5329 7644
rect 5353 7642 5409 7644
rect 5433 7642 5489 7644
rect 5513 7642 5569 7644
rect 5273 7590 5319 7642
rect 5319 7590 5329 7642
rect 5353 7590 5383 7642
rect 5383 7590 5395 7642
rect 5395 7590 5409 7642
rect 5433 7590 5447 7642
rect 5447 7590 5459 7642
rect 5459 7590 5489 7642
rect 5513 7590 5523 7642
rect 5523 7590 5569 7642
rect 5273 7588 5329 7590
rect 5353 7588 5409 7590
rect 5433 7588 5489 7590
rect 5513 7588 5569 7590
rect 4613 7098 4669 7100
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4613 7046 4659 7098
rect 4659 7046 4669 7098
rect 4693 7046 4723 7098
rect 4723 7046 4735 7098
rect 4735 7046 4749 7098
rect 4773 7046 4787 7098
rect 4787 7046 4799 7098
rect 4799 7046 4829 7098
rect 4853 7046 4863 7098
rect 4863 7046 4909 7098
rect 4613 7044 4669 7046
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 5273 6554 5329 6556
rect 5353 6554 5409 6556
rect 5433 6554 5489 6556
rect 5513 6554 5569 6556
rect 5273 6502 5319 6554
rect 5319 6502 5329 6554
rect 5353 6502 5383 6554
rect 5383 6502 5395 6554
rect 5395 6502 5409 6554
rect 5433 6502 5447 6554
rect 5447 6502 5459 6554
rect 5459 6502 5489 6554
rect 5513 6502 5523 6554
rect 5523 6502 5569 6554
rect 5273 6500 5329 6502
rect 5353 6500 5409 6502
rect 5433 6500 5489 6502
rect 5513 6500 5569 6502
rect 4613 6010 4669 6012
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4613 5958 4659 6010
rect 4659 5958 4669 6010
rect 4693 5958 4723 6010
rect 4723 5958 4735 6010
rect 4735 5958 4749 6010
rect 4773 5958 4787 6010
rect 4787 5958 4799 6010
rect 4799 5958 4829 6010
rect 4853 5958 4863 6010
rect 4863 5958 4909 6010
rect 4613 5956 4669 5958
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4613 4922 4669 4924
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4613 4870 4659 4922
rect 4659 4870 4669 4922
rect 4693 4870 4723 4922
rect 4723 4870 4735 4922
rect 4735 4870 4749 4922
rect 4773 4870 4787 4922
rect 4787 4870 4799 4922
rect 4799 4870 4829 4922
rect 4853 4870 4863 4922
rect 4863 4870 4909 4922
rect 4613 4868 4669 4870
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 2835 4378 2891 4380
rect 2915 4378 2971 4380
rect 2995 4378 3051 4380
rect 3075 4378 3131 4380
rect 2835 4326 2881 4378
rect 2881 4326 2891 4378
rect 2915 4326 2945 4378
rect 2945 4326 2957 4378
rect 2957 4326 2971 4378
rect 2995 4326 3009 4378
rect 3009 4326 3021 4378
rect 3021 4326 3051 4378
rect 3075 4326 3085 4378
rect 3085 4326 3131 4378
rect 2835 4324 2891 4326
rect 2915 4324 2971 4326
rect 2995 4324 3051 4326
rect 3075 4324 3131 4326
rect 846 3576 848 3596
rect 848 3576 900 3596
rect 900 3576 902 3596
rect 2594 3576 2650 3632
rect 5273 5466 5329 5468
rect 5353 5466 5409 5468
rect 5433 5466 5489 5468
rect 5513 5466 5569 5468
rect 5273 5414 5319 5466
rect 5319 5414 5329 5466
rect 5353 5414 5383 5466
rect 5383 5414 5395 5466
rect 5395 5414 5409 5466
rect 5433 5414 5447 5466
rect 5447 5414 5459 5466
rect 5459 5414 5489 5466
rect 5513 5414 5523 5466
rect 5523 5414 5569 5466
rect 5273 5412 5329 5414
rect 5353 5412 5409 5414
rect 5433 5412 5489 5414
rect 5513 5412 5569 5414
rect 5273 4378 5329 4380
rect 5353 4378 5409 4380
rect 5433 4378 5489 4380
rect 5513 4378 5569 4380
rect 5273 4326 5319 4378
rect 5319 4326 5329 4378
rect 5353 4326 5383 4378
rect 5383 4326 5395 4378
rect 5395 4326 5409 4378
rect 5433 4326 5447 4378
rect 5447 4326 5459 4378
rect 5459 4326 5489 4378
rect 5513 4326 5523 4378
rect 5523 4326 5569 4378
rect 5273 4324 5329 4326
rect 5353 4324 5409 4326
rect 5433 4324 5489 4326
rect 5513 4324 5569 4326
rect 7051 10362 7107 10364
rect 7131 10362 7187 10364
rect 7211 10362 7267 10364
rect 7291 10362 7347 10364
rect 7051 10310 7097 10362
rect 7097 10310 7107 10362
rect 7131 10310 7161 10362
rect 7161 10310 7173 10362
rect 7173 10310 7187 10362
rect 7211 10310 7225 10362
rect 7225 10310 7237 10362
rect 7237 10310 7267 10362
rect 7291 10310 7301 10362
rect 7301 10310 7347 10362
rect 7051 10308 7107 10310
rect 7131 10308 7187 10310
rect 7211 10308 7267 10310
rect 7291 10308 7347 10310
rect 9489 11450 9545 11452
rect 9569 11450 9625 11452
rect 9649 11450 9705 11452
rect 9729 11450 9785 11452
rect 9489 11398 9535 11450
rect 9535 11398 9545 11450
rect 9569 11398 9599 11450
rect 9599 11398 9611 11450
rect 9611 11398 9625 11450
rect 9649 11398 9663 11450
rect 9663 11398 9675 11450
rect 9675 11398 9705 11450
rect 9729 11398 9739 11450
rect 9739 11398 9785 11450
rect 9489 11396 9545 11398
rect 9569 11396 9625 11398
rect 9649 11396 9705 11398
rect 9729 11396 9785 11398
rect 10149 10906 10205 10908
rect 10229 10906 10285 10908
rect 10309 10906 10365 10908
rect 10389 10906 10445 10908
rect 10149 10854 10195 10906
rect 10195 10854 10205 10906
rect 10229 10854 10259 10906
rect 10259 10854 10271 10906
rect 10271 10854 10285 10906
rect 10309 10854 10323 10906
rect 10323 10854 10335 10906
rect 10335 10854 10365 10906
rect 10389 10854 10399 10906
rect 10399 10854 10445 10906
rect 10149 10852 10205 10854
rect 10229 10852 10285 10854
rect 10309 10852 10365 10854
rect 10389 10852 10445 10854
rect 7711 9818 7767 9820
rect 7791 9818 7847 9820
rect 7871 9818 7927 9820
rect 7951 9818 8007 9820
rect 7711 9766 7757 9818
rect 7757 9766 7767 9818
rect 7791 9766 7821 9818
rect 7821 9766 7833 9818
rect 7833 9766 7847 9818
rect 7871 9766 7885 9818
rect 7885 9766 7897 9818
rect 7897 9766 7927 9818
rect 7951 9766 7961 9818
rect 7961 9766 8007 9818
rect 7711 9764 7767 9766
rect 7791 9764 7847 9766
rect 7871 9764 7927 9766
rect 7951 9764 8007 9766
rect 9489 10362 9545 10364
rect 9569 10362 9625 10364
rect 9649 10362 9705 10364
rect 9729 10362 9785 10364
rect 9489 10310 9535 10362
rect 9535 10310 9545 10362
rect 9569 10310 9599 10362
rect 9599 10310 9611 10362
rect 9611 10310 9625 10362
rect 9649 10310 9663 10362
rect 9663 10310 9675 10362
rect 9675 10310 9705 10362
rect 9729 10310 9739 10362
rect 9739 10310 9785 10362
rect 9489 10308 9545 10310
rect 9569 10308 9625 10310
rect 9649 10308 9705 10310
rect 9729 10308 9785 10310
rect 10149 9818 10205 9820
rect 10229 9818 10285 9820
rect 10309 9818 10365 9820
rect 10389 9818 10445 9820
rect 10149 9766 10195 9818
rect 10195 9766 10205 9818
rect 10229 9766 10259 9818
rect 10259 9766 10271 9818
rect 10271 9766 10285 9818
rect 10309 9766 10323 9818
rect 10323 9766 10335 9818
rect 10335 9766 10365 9818
rect 10389 9766 10399 9818
rect 10399 9766 10445 9818
rect 10149 9764 10205 9766
rect 10229 9764 10285 9766
rect 10309 9764 10365 9766
rect 10389 9764 10445 9766
rect 7051 9274 7107 9276
rect 7131 9274 7187 9276
rect 7211 9274 7267 9276
rect 7291 9274 7347 9276
rect 7051 9222 7097 9274
rect 7097 9222 7107 9274
rect 7131 9222 7161 9274
rect 7161 9222 7173 9274
rect 7173 9222 7187 9274
rect 7211 9222 7225 9274
rect 7225 9222 7237 9274
rect 7237 9222 7267 9274
rect 7291 9222 7301 9274
rect 7301 9222 7347 9274
rect 7051 9220 7107 9222
rect 7131 9220 7187 9222
rect 7211 9220 7267 9222
rect 7291 9220 7347 9222
rect 7051 8186 7107 8188
rect 7131 8186 7187 8188
rect 7211 8186 7267 8188
rect 7291 8186 7347 8188
rect 7051 8134 7097 8186
rect 7097 8134 7107 8186
rect 7131 8134 7161 8186
rect 7161 8134 7173 8186
rect 7173 8134 7187 8186
rect 7211 8134 7225 8186
rect 7225 8134 7237 8186
rect 7237 8134 7267 8186
rect 7291 8134 7301 8186
rect 7301 8134 7347 8186
rect 7051 8132 7107 8134
rect 7131 8132 7187 8134
rect 7211 8132 7267 8134
rect 7291 8132 7347 8134
rect 9489 9274 9545 9276
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9489 9222 9535 9274
rect 9535 9222 9545 9274
rect 9569 9222 9599 9274
rect 9599 9222 9611 9274
rect 9611 9222 9625 9274
rect 9649 9222 9663 9274
rect 9663 9222 9675 9274
rect 9675 9222 9705 9274
rect 9729 9222 9739 9274
rect 9739 9222 9785 9274
rect 9489 9220 9545 9222
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 10506 8916 10508 8936
rect 10508 8916 10560 8936
rect 10560 8916 10562 8936
rect 7711 8730 7767 8732
rect 7791 8730 7847 8732
rect 7871 8730 7927 8732
rect 7951 8730 8007 8732
rect 7711 8678 7757 8730
rect 7757 8678 7767 8730
rect 7791 8678 7821 8730
rect 7821 8678 7833 8730
rect 7833 8678 7847 8730
rect 7871 8678 7885 8730
rect 7885 8678 7897 8730
rect 7897 8678 7927 8730
rect 7951 8678 7961 8730
rect 7961 8678 8007 8730
rect 7711 8676 7767 8678
rect 7791 8676 7847 8678
rect 7871 8676 7927 8678
rect 7951 8676 8007 8678
rect 7711 7642 7767 7644
rect 7791 7642 7847 7644
rect 7871 7642 7927 7644
rect 7951 7642 8007 7644
rect 7711 7590 7757 7642
rect 7757 7590 7767 7642
rect 7791 7590 7821 7642
rect 7821 7590 7833 7642
rect 7833 7590 7847 7642
rect 7871 7590 7885 7642
rect 7885 7590 7897 7642
rect 7897 7590 7927 7642
rect 7951 7590 7961 7642
rect 7961 7590 8007 7642
rect 7711 7588 7767 7590
rect 7791 7588 7847 7590
rect 7871 7588 7927 7590
rect 7951 7588 8007 7590
rect 7051 7098 7107 7100
rect 7131 7098 7187 7100
rect 7211 7098 7267 7100
rect 7291 7098 7347 7100
rect 7051 7046 7097 7098
rect 7097 7046 7107 7098
rect 7131 7046 7161 7098
rect 7161 7046 7173 7098
rect 7173 7046 7187 7098
rect 7211 7046 7225 7098
rect 7225 7046 7237 7098
rect 7237 7046 7267 7098
rect 7291 7046 7301 7098
rect 7301 7046 7347 7098
rect 7051 7044 7107 7046
rect 7131 7044 7187 7046
rect 7211 7044 7267 7046
rect 7291 7044 7347 7046
rect 7051 6010 7107 6012
rect 7131 6010 7187 6012
rect 7211 6010 7267 6012
rect 7291 6010 7347 6012
rect 7051 5958 7097 6010
rect 7097 5958 7107 6010
rect 7131 5958 7161 6010
rect 7161 5958 7173 6010
rect 7173 5958 7187 6010
rect 7211 5958 7225 6010
rect 7225 5958 7237 6010
rect 7237 5958 7267 6010
rect 7291 5958 7301 6010
rect 7301 5958 7347 6010
rect 7051 5956 7107 5958
rect 7131 5956 7187 5958
rect 7211 5956 7267 5958
rect 7291 5956 7347 5958
rect 6826 5208 6882 5264
rect 3514 3596 3570 3632
rect 3514 3576 3516 3596
rect 3516 3576 3568 3596
rect 3568 3576 3570 3596
rect 2835 3290 2891 3292
rect 2915 3290 2971 3292
rect 2995 3290 3051 3292
rect 3075 3290 3131 3292
rect 2835 3238 2881 3290
rect 2881 3238 2891 3290
rect 2915 3238 2945 3290
rect 2945 3238 2957 3290
rect 2957 3238 2971 3290
rect 2995 3238 3009 3290
rect 3009 3238 3021 3290
rect 3021 3238 3051 3290
rect 3075 3238 3085 3290
rect 3085 3238 3131 3290
rect 2835 3236 2891 3238
rect 2915 3236 2971 3238
rect 2995 3236 3051 3238
rect 3075 3236 3131 3238
rect 4066 3052 4122 3088
rect 4066 3032 4068 3052
rect 4068 3032 4120 3052
rect 4120 3032 4122 3052
rect 4613 3834 4669 3836
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4613 3782 4659 3834
rect 4659 3782 4669 3834
rect 4693 3782 4723 3834
rect 4723 3782 4735 3834
rect 4735 3782 4749 3834
rect 4773 3782 4787 3834
rect 4787 3782 4799 3834
rect 4799 3782 4829 3834
rect 4853 3782 4863 3834
rect 4863 3782 4909 3834
rect 4613 3780 4669 3782
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 2175 2746 2231 2748
rect 2255 2746 2311 2748
rect 2335 2746 2391 2748
rect 2415 2746 2471 2748
rect 2175 2694 2221 2746
rect 2221 2694 2231 2746
rect 2255 2694 2285 2746
rect 2285 2694 2297 2746
rect 2297 2694 2311 2746
rect 2335 2694 2349 2746
rect 2349 2694 2361 2746
rect 2361 2694 2391 2746
rect 2415 2694 2425 2746
rect 2425 2694 2471 2746
rect 2175 2692 2231 2694
rect 2255 2692 2311 2694
rect 2335 2692 2391 2694
rect 2415 2692 2471 2694
rect 5273 3290 5329 3292
rect 5353 3290 5409 3292
rect 5433 3290 5489 3292
rect 5513 3290 5569 3292
rect 5273 3238 5319 3290
rect 5319 3238 5329 3290
rect 5353 3238 5383 3290
rect 5383 3238 5395 3290
rect 5395 3238 5409 3290
rect 5433 3238 5447 3290
rect 5447 3238 5459 3290
rect 5459 3238 5489 3290
rect 5513 3238 5523 3290
rect 5523 3238 5569 3290
rect 5273 3236 5329 3238
rect 5353 3236 5409 3238
rect 5433 3236 5489 3238
rect 5513 3236 5569 3238
rect 4613 2746 4669 2748
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4613 2694 4659 2746
rect 4659 2694 4669 2746
rect 4693 2694 4723 2746
rect 4723 2694 4735 2746
rect 4735 2694 4749 2746
rect 4773 2694 4787 2746
rect 4787 2694 4799 2746
rect 4799 2694 4829 2746
rect 4853 2694 4863 2746
rect 4863 2694 4909 2746
rect 4613 2692 4669 2694
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 7051 4922 7107 4924
rect 7131 4922 7187 4924
rect 7211 4922 7267 4924
rect 7291 4922 7347 4924
rect 7051 4870 7097 4922
rect 7097 4870 7107 4922
rect 7131 4870 7161 4922
rect 7161 4870 7173 4922
rect 7173 4870 7187 4922
rect 7211 4870 7225 4922
rect 7225 4870 7237 4922
rect 7237 4870 7267 4922
rect 7291 4870 7301 4922
rect 7301 4870 7347 4922
rect 7051 4868 7107 4870
rect 7131 4868 7187 4870
rect 7211 4868 7267 4870
rect 7291 4868 7347 4870
rect 7711 6554 7767 6556
rect 7791 6554 7847 6556
rect 7871 6554 7927 6556
rect 7951 6554 8007 6556
rect 7711 6502 7757 6554
rect 7757 6502 7767 6554
rect 7791 6502 7821 6554
rect 7821 6502 7833 6554
rect 7833 6502 7847 6554
rect 7871 6502 7885 6554
rect 7885 6502 7897 6554
rect 7897 6502 7927 6554
rect 7951 6502 7961 6554
rect 7961 6502 8007 6554
rect 7711 6500 7767 6502
rect 7791 6500 7847 6502
rect 7871 6500 7927 6502
rect 7951 6500 8007 6502
rect 7470 5228 7526 5264
rect 7470 5208 7472 5228
rect 7472 5208 7524 5228
rect 7524 5208 7526 5228
rect 7051 3834 7107 3836
rect 7131 3834 7187 3836
rect 7211 3834 7267 3836
rect 7291 3834 7347 3836
rect 7051 3782 7097 3834
rect 7097 3782 7107 3834
rect 7131 3782 7161 3834
rect 7161 3782 7173 3834
rect 7173 3782 7187 3834
rect 7211 3782 7225 3834
rect 7225 3782 7237 3834
rect 7237 3782 7267 3834
rect 7291 3782 7301 3834
rect 7301 3782 7347 3834
rect 7051 3780 7107 3782
rect 7131 3780 7187 3782
rect 7211 3780 7267 3782
rect 7291 3780 7347 3782
rect 7711 5466 7767 5468
rect 7791 5466 7847 5468
rect 7871 5466 7927 5468
rect 7951 5466 8007 5468
rect 7711 5414 7757 5466
rect 7757 5414 7767 5466
rect 7791 5414 7821 5466
rect 7821 5414 7833 5466
rect 7833 5414 7847 5466
rect 7871 5414 7885 5466
rect 7885 5414 7897 5466
rect 7897 5414 7927 5466
rect 7951 5414 7961 5466
rect 7961 5414 8007 5466
rect 7711 5412 7767 5414
rect 7791 5412 7847 5414
rect 7871 5412 7927 5414
rect 7951 5412 8007 5414
rect 7470 3576 7526 3632
rect 10506 8880 10562 8916
rect 10149 8730 10205 8732
rect 10229 8730 10285 8732
rect 10309 8730 10365 8732
rect 10389 8730 10445 8732
rect 10149 8678 10195 8730
rect 10195 8678 10205 8730
rect 10229 8678 10259 8730
rect 10259 8678 10271 8730
rect 10271 8678 10285 8730
rect 10309 8678 10323 8730
rect 10323 8678 10335 8730
rect 10335 8678 10365 8730
rect 10389 8678 10399 8730
rect 10399 8678 10445 8730
rect 10149 8676 10205 8678
rect 10229 8676 10285 8678
rect 10309 8676 10365 8678
rect 10389 8676 10445 8678
rect 9489 8186 9545 8188
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9489 8134 9535 8186
rect 9535 8134 9545 8186
rect 9569 8134 9599 8186
rect 9599 8134 9611 8186
rect 9611 8134 9625 8186
rect 9649 8134 9663 8186
rect 9663 8134 9675 8186
rect 9675 8134 9705 8186
rect 9729 8134 9739 8186
rect 9739 8134 9785 8186
rect 9489 8132 9545 8134
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 10506 8200 10562 8256
rect 9489 7098 9545 7100
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9489 7046 9535 7098
rect 9535 7046 9545 7098
rect 9569 7046 9599 7098
rect 9599 7046 9611 7098
rect 9611 7046 9625 7098
rect 9649 7046 9663 7098
rect 9663 7046 9675 7098
rect 9675 7046 9705 7098
rect 9729 7046 9739 7098
rect 9739 7046 9785 7098
rect 9489 7044 9545 7046
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 10149 7642 10205 7644
rect 10229 7642 10285 7644
rect 10309 7642 10365 7644
rect 10389 7642 10445 7644
rect 10149 7590 10195 7642
rect 10195 7590 10205 7642
rect 10229 7590 10259 7642
rect 10259 7590 10271 7642
rect 10271 7590 10285 7642
rect 10309 7590 10323 7642
rect 10323 7590 10335 7642
rect 10335 7590 10365 7642
rect 10389 7590 10399 7642
rect 10399 7590 10445 7642
rect 10149 7588 10205 7590
rect 10229 7588 10285 7590
rect 10309 7588 10365 7590
rect 10389 7588 10445 7590
rect 10690 7520 10746 7576
rect 10414 6840 10470 6896
rect 7711 4378 7767 4380
rect 7791 4378 7847 4380
rect 7871 4378 7927 4380
rect 7951 4378 8007 4380
rect 7711 4326 7757 4378
rect 7757 4326 7767 4378
rect 7791 4326 7821 4378
rect 7821 4326 7833 4378
rect 7833 4326 7847 4378
rect 7871 4326 7885 4378
rect 7885 4326 7897 4378
rect 7897 4326 7927 4378
rect 7951 4326 7961 4378
rect 7961 4326 8007 4378
rect 7711 4324 7767 4326
rect 7791 4324 7847 4326
rect 7871 4324 7927 4326
rect 7951 4324 8007 4326
rect 9489 6010 9545 6012
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9489 5958 9535 6010
rect 9535 5958 9545 6010
rect 9569 5958 9599 6010
rect 9599 5958 9611 6010
rect 9611 5958 9625 6010
rect 9649 5958 9663 6010
rect 9663 5958 9675 6010
rect 9675 5958 9705 6010
rect 9729 5958 9739 6010
rect 9739 5958 9785 6010
rect 9489 5956 9545 5958
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 10149 6554 10205 6556
rect 10229 6554 10285 6556
rect 10309 6554 10365 6556
rect 10389 6554 10445 6556
rect 10149 6502 10195 6554
rect 10195 6502 10205 6554
rect 10229 6502 10259 6554
rect 10259 6502 10271 6554
rect 10271 6502 10285 6554
rect 10309 6502 10323 6554
rect 10323 6502 10335 6554
rect 10335 6502 10365 6554
rect 10389 6502 10399 6554
rect 10399 6502 10445 6554
rect 10149 6500 10205 6502
rect 10229 6500 10285 6502
rect 10309 6500 10365 6502
rect 10389 6500 10445 6502
rect 9489 4922 9545 4924
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9489 4870 9535 4922
rect 9535 4870 9545 4922
rect 9569 4870 9599 4922
rect 9599 4870 9611 4922
rect 9611 4870 9625 4922
rect 9649 4870 9663 4922
rect 9663 4870 9675 4922
rect 9675 4870 9705 4922
rect 9729 4870 9739 4922
rect 9739 4870 9785 4922
rect 9489 4868 9545 4870
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 7102 3032 7158 3088
rect 7711 3290 7767 3292
rect 7791 3290 7847 3292
rect 7871 3290 7927 3292
rect 7951 3290 8007 3292
rect 7711 3238 7757 3290
rect 7757 3238 7767 3290
rect 7791 3238 7821 3290
rect 7821 3238 7833 3290
rect 7833 3238 7847 3290
rect 7871 3238 7885 3290
rect 7885 3238 7897 3290
rect 7897 3238 7927 3290
rect 7951 3238 7961 3290
rect 7961 3238 8007 3290
rect 7711 3236 7767 3238
rect 7791 3236 7847 3238
rect 7871 3236 7927 3238
rect 7951 3236 8007 3238
rect 9489 3834 9545 3836
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9489 3782 9535 3834
rect 9535 3782 9545 3834
rect 9569 3782 9599 3834
rect 9599 3782 9611 3834
rect 9611 3782 9625 3834
rect 9649 3782 9663 3834
rect 9663 3782 9675 3834
rect 9675 3782 9705 3834
rect 9729 3782 9739 3834
rect 9739 3782 9785 3834
rect 9489 3780 9545 3782
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 7051 2746 7107 2748
rect 7131 2746 7187 2748
rect 7211 2746 7267 2748
rect 7291 2746 7347 2748
rect 7051 2694 7097 2746
rect 7097 2694 7107 2746
rect 7131 2694 7161 2746
rect 7161 2694 7173 2746
rect 7173 2694 7187 2746
rect 7211 2694 7225 2746
rect 7225 2694 7237 2746
rect 7237 2694 7267 2746
rect 7291 2694 7301 2746
rect 7301 2694 7347 2746
rect 7051 2692 7107 2694
rect 7131 2692 7187 2694
rect 7211 2692 7267 2694
rect 7291 2692 7347 2694
rect 10414 6160 10470 6216
rect 10598 5480 10654 5536
rect 10149 5466 10205 5468
rect 10229 5466 10285 5468
rect 10309 5466 10365 5468
rect 10389 5466 10445 5468
rect 10149 5414 10195 5466
rect 10195 5414 10205 5466
rect 10229 5414 10259 5466
rect 10259 5414 10271 5466
rect 10271 5414 10285 5466
rect 10309 5414 10323 5466
rect 10323 5414 10335 5466
rect 10335 5414 10365 5466
rect 10389 5414 10399 5466
rect 10399 5414 10445 5466
rect 10149 5412 10205 5414
rect 10229 5412 10285 5414
rect 10309 5412 10365 5414
rect 10389 5412 10445 5414
rect 10506 4800 10562 4856
rect 10149 4378 10205 4380
rect 10229 4378 10285 4380
rect 10309 4378 10365 4380
rect 10389 4378 10445 4380
rect 10149 4326 10195 4378
rect 10195 4326 10205 4378
rect 10229 4326 10259 4378
rect 10259 4326 10271 4378
rect 10271 4326 10285 4378
rect 10309 4326 10323 4378
rect 10323 4326 10335 4378
rect 10335 4326 10365 4378
rect 10389 4326 10399 4378
rect 10399 4326 10445 4378
rect 10149 4324 10205 4326
rect 10229 4324 10285 4326
rect 10309 4324 10365 4326
rect 10389 4324 10445 4326
rect 10149 3290 10205 3292
rect 10229 3290 10285 3292
rect 10309 3290 10365 3292
rect 10389 3290 10445 3292
rect 10149 3238 10195 3290
rect 10195 3238 10205 3290
rect 10229 3238 10259 3290
rect 10259 3238 10271 3290
rect 10271 3238 10285 3290
rect 10309 3238 10323 3290
rect 10323 3238 10335 3290
rect 10335 3238 10365 3290
rect 10389 3238 10399 3290
rect 10399 3238 10445 3290
rect 10149 3236 10205 3238
rect 10229 3236 10285 3238
rect 10309 3236 10365 3238
rect 10389 3236 10445 3238
rect 9489 2746 9545 2748
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9489 2694 9535 2746
rect 9535 2694 9545 2746
rect 9569 2694 9599 2746
rect 9599 2694 9611 2746
rect 9611 2694 9625 2746
rect 9649 2694 9663 2746
rect 9663 2694 9675 2746
rect 9675 2694 9705 2746
rect 9729 2694 9739 2746
rect 9739 2694 9785 2746
rect 9489 2692 9545 2694
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 2835 2202 2891 2204
rect 2915 2202 2971 2204
rect 2995 2202 3051 2204
rect 3075 2202 3131 2204
rect 2835 2150 2881 2202
rect 2881 2150 2891 2202
rect 2915 2150 2945 2202
rect 2945 2150 2957 2202
rect 2957 2150 2971 2202
rect 2995 2150 3009 2202
rect 3009 2150 3021 2202
rect 3021 2150 3051 2202
rect 3075 2150 3085 2202
rect 3085 2150 3131 2202
rect 2835 2148 2891 2150
rect 2915 2148 2971 2150
rect 2995 2148 3051 2150
rect 3075 2148 3131 2150
rect 5273 2202 5329 2204
rect 5353 2202 5409 2204
rect 5433 2202 5489 2204
rect 5513 2202 5569 2204
rect 5273 2150 5319 2202
rect 5319 2150 5329 2202
rect 5353 2150 5383 2202
rect 5383 2150 5395 2202
rect 5395 2150 5409 2202
rect 5433 2150 5447 2202
rect 5447 2150 5459 2202
rect 5459 2150 5489 2202
rect 5513 2150 5523 2202
rect 5523 2150 5569 2202
rect 5273 2148 5329 2150
rect 5353 2148 5409 2150
rect 5433 2148 5489 2150
rect 5513 2148 5569 2150
rect 7711 2202 7767 2204
rect 7791 2202 7847 2204
rect 7871 2202 7927 2204
rect 7951 2202 8007 2204
rect 7711 2150 7757 2202
rect 7757 2150 7767 2202
rect 7791 2150 7821 2202
rect 7821 2150 7833 2202
rect 7833 2150 7847 2202
rect 7871 2150 7885 2202
rect 7885 2150 7897 2202
rect 7897 2150 7927 2202
rect 7951 2150 7961 2202
rect 7961 2150 8007 2202
rect 7711 2148 7767 2150
rect 7791 2148 7847 2150
rect 7871 2148 7927 2150
rect 7951 2148 8007 2150
rect 10149 2202 10205 2204
rect 10229 2202 10285 2204
rect 10309 2202 10365 2204
rect 10389 2202 10445 2204
rect 10149 2150 10195 2202
rect 10195 2150 10205 2202
rect 10229 2150 10259 2202
rect 10259 2150 10271 2202
rect 10271 2150 10285 2202
rect 10309 2150 10323 2202
rect 10323 2150 10335 2202
rect 10335 2150 10365 2202
rect 10389 2150 10399 2202
rect 10399 2150 10445 2202
rect 10149 2148 10205 2150
rect 10229 2148 10285 2150
rect 10309 2148 10365 2150
rect 10389 2148 10445 2150
<< metal3 >>
rect 2165 11456 2481 11457
rect 2165 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2481 11456
rect 2165 11391 2481 11392
rect 4603 11456 4919 11457
rect 4603 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4919 11456
rect 4603 11391 4919 11392
rect 7041 11456 7357 11457
rect 7041 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7357 11456
rect 7041 11391 7357 11392
rect 9479 11456 9795 11457
rect 9479 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9795 11456
rect 9479 11391 9795 11392
rect 2825 10912 3141 10913
rect 2825 10848 2831 10912
rect 2895 10848 2911 10912
rect 2975 10848 2991 10912
rect 3055 10848 3071 10912
rect 3135 10848 3141 10912
rect 2825 10847 3141 10848
rect 5263 10912 5579 10913
rect 5263 10848 5269 10912
rect 5333 10848 5349 10912
rect 5413 10848 5429 10912
rect 5493 10848 5509 10912
rect 5573 10848 5579 10912
rect 5263 10847 5579 10848
rect 7701 10912 8017 10913
rect 7701 10848 7707 10912
rect 7771 10848 7787 10912
rect 7851 10848 7867 10912
rect 7931 10848 7947 10912
rect 8011 10848 8017 10912
rect 7701 10847 8017 10848
rect 10139 10912 10455 10913
rect 10139 10848 10145 10912
rect 10209 10848 10225 10912
rect 10289 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10455 10912
rect 10139 10847 10455 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 2165 10368 2481 10369
rect 2165 10304 2171 10368
rect 2235 10304 2251 10368
rect 2315 10304 2331 10368
rect 2395 10304 2411 10368
rect 2475 10304 2481 10368
rect 2165 10303 2481 10304
rect 4603 10368 4919 10369
rect 4603 10304 4609 10368
rect 4673 10304 4689 10368
rect 4753 10304 4769 10368
rect 4833 10304 4849 10368
rect 4913 10304 4919 10368
rect 4603 10303 4919 10304
rect 7041 10368 7357 10369
rect 7041 10304 7047 10368
rect 7111 10304 7127 10368
rect 7191 10304 7207 10368
rect 7271 10304 7287 10368
rect 7351 10304 7357 10368
rect 7041 10303 7357 10304
rect 9479 10368 9795 10369
rect 9479 10304 9485 10368
rect 9549 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9795 10368
rect 9479 10303 9795 10304
rect 0 10208 800 10238
rect 2825 9824 3141 9825
rect 2825 9760 2831 9824
rect 2895 9760 2911 9824
rect 2975 9760 2991 9824
rect 3055 9760 3071 9824
rect 3135 9760 3141 9824
rect 2825 9759 3141 9760
rect 5263 9824 5579 9825
rect 5263 9760 5269 9824
rect 5333 9760 5349 9824
rect 5413 9760 5429 9824
rect 5493 9760 5509 9824
rect 5573 9760 5579 9824
rect 5263 9759 5579 9760
rect 7701 9824 8017 9825
rect 7701 9760 7707 9824
rect 7771 9760 7787 9824
rect 7851 9760 7867 9824
rect 7931 9760 7947 9824
rect 8011 9760 8017 9824
rect 7701 9759 8017 9760
rect 10139 9824 10455 9825
rect 10139 9760 10145 9824
rect 10209 9760 10225 9824
rect 10289 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10455 9824
rect 10139 9759 10455 9760
rect 2165 9280 2481 9281
rect 2165 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2481 9280
rect 2165 9215 2481 9216
rect 4603 9280 4919 9281
rect 4603 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4919 9280
rect 4603 9215 4919 9216
rect 7041 9280 7357 9281
rect 7041 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7357 9280
rect 7041 9215 7357 9216
rect 9479 9280 9795 9281
rect 9479 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9795 9280
rect 9479 9215 9795 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 10501 8938 10567 8941
rect 11198 8938 11998 8968
rect 10501 8936 11998 8938
rect 10501 8880 10506 8936
rect 10562 8880 11998 8936
rect 10501 8878 11998 8880
rect 0 8848 800 8878
rect 10501 8875 10567 8878
rect 11198 8848 11998 8878
rect 2825 8736 3141 8737
rect 2825 8672 2831 8736
rect 2895 8672 2911 8736
rect 2975 8672 2991 8736
rect 3055 8672 3071 8736
rect 3135 8672 3141 8736
rect 2825 8671 3141 8672
rect 5263 8736 5579 8737
rect 5263 8672 5269 8736
rect 5333 8672 5349 8736
rect 5413 8672 5429 8736
rect 5493 8672 5509 8736
rect 5573 8672 5579 8736
rect 5263 8671 5579 8672
rect 7701 8736 8017 8737
rect 7701 8672 7707 8736
rect 7771 8672 7787 8736
rect 7851 8672 7867 8736
rect 7931 8672 7947 8736
rect 8011 8672 8017 8736
rect 7701 8671 8017 8672
rect 10139 8736 10455 8737
rect 10139 8672 10145 8736
rect 10209 8672 10225 8736
rect 10289 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10455 8736
rect 10139 8671 10455 8672
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 10501 8258 10567 8261
rect 11198 8258 11998 8288
rect 10501 8256 11998 8258
rect 10501 8200 10506 8256
rect 10562 8200 11998 8256
rect 10501 8198 11998 8200
rect 10501 8195 10567 8198
rect 2165 8192 2481 8193
rect 2165 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2481 8192
rect 2165 8127 2481 8128
rect 4603 8192 4919 8193
rect 4603 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4919 8192
rect 4603 8127 4919 8128
rect 7041 8192 7357 8193
rect 7041 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7357 8192
rect 7041 8127 7357 8128
rect 9479 8192 9795 8193
rect 9479 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9795 8192
rect 11198 8168 11998 8198
rect 9479 8127 9795 8128
rect 2825 7648 3141 7649
rect 0 7578 800 7608
rect 2825 7584 2831 7648
rect 2895 7584 2911 7648
rect 2975 7584 2991 7648
rect 3055 7584 3071 7648
rect 3135 7584 3141 7648
rect 2825 7583 3141 7584
rect 5263 7648 5579 7649
rect 5263 7584 5269 7648
rect 5333 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5579 7648
rect 5263 7583 5579 7584
rect 7701 7648 8017 7649
rect 7701 7584 7707 7648
rect 7771 7584 7787 7648
rect 7851 7584 7867 7648
rect 7931 7584 7947 7648
rect 8011 7584 8017 7648
rect 7701 7583 8017 7584
rect 10139 7648 10455 7649
rect 10139 7584 10145 7648
rect 10209 7584 10225 7648
rect 10289 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10455 7648
rect 10139 7583 10455 7584
rect 10685 7578 10751 7581
rect 11198 7578 11998 7608
rect 0 7488 858 7578
rect 10685 7576 11998 7578
rect 10685 7520 10690 7576
rect 10746 7520 11998 7576
rect 10685 7518 11998 7520
rect 10685 7515 10751 7518
rect 11198 7488 11998 7518
rect 798 7445 858 7488
rect 798 7440 907 7445
rect 798 7384 846 7440
rect 902 7384 907 7440
rect 798 7382 907 7384
rect 841 7379 907 7382
rect 2165 7104 2481 7105
rect 2165 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2481 7104
rect 2165 7039 2481 7040
rect 4603 7104 4919 7105
rect 4603 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4919 7104
rect 4603 7039 4919 7040
rect 7041 7104 7357 7105
rect 7041 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7357 7104
rect 7041 7039 7357 7040
rect 9479 7104 9795 7105
rect 9479 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9795 7104
rect 9479 7039 9795 7040
rect 10409 6898 10475 6901
rect 11198 6898 11998 6928
rect 10409 6896 11998 6898
rect 10409 6840 10414 6896
rect 10470 6840 11998 6896
rect 10409 6838 11998 6840
rect 10409 6835 10475 6838
rect 11198 6808 11998 6838
rect 2825 6560 3141 6561
rect 2825 6496 2831 6560
rect 2895 6496 2911 6560
rect 2975 6496 2991 6560
rect 3055 6496 3071 6560
rect 3135 6496 3141 6560
rect 2825 6495 3141 6496
rect 5263 6560 5579 6561
rect 5263 6496 5269 6560
rect 5333 6496 5349 6560
rect 5413 6496 5429 6560
rect 5493 6496 5509 6560
rect 5573 6496 5579 6560
rect 5263 6495 5579 6496
rect 7701 6560 8017 6561
rect 7701 6496 7707 6560
rect 7771 6496 7787 6560
rect 7851 6496 7867 6560
rect 7931 6496 7947 6560
rect 8011 6496 8017 6560
rect 7701 6495 8017 6496
rect 10139 6560 10455 6561
rect 10139 6496 10145 6560
rect 10209 6496 10225 6560
rect 10289 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10455 6560
rect 10139 6495 10455 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 10409 6218 10475 6221
rect 11198 6218 11998 6248
rect 10409 6216 11998 6218
rect 10409 6160 10414 6216
rect 10470 6160 11998 6216
rect 10409 6158 11998 6160
rect 0 6128 800 6158
rect 10409 6155 10475 6158
rect 11198 6128 11998 6158
rect 2165 6016 2481 6017
rect 2165 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2481 6016
rect 2165 5951 2481 5952
rect 4603 6016 4919 6017
rect 4603 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4919 6016
rect 4603 5951 4919 5952
rect 7041 6016 7357 6017
rect 7041 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7357 6016
rect 7041 5951 7357 5952
rect 9479 6016 9795 6017
rect 9479 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9795 6016
rect 9479 5951 9795 5952
rect 0 5538 800 5568
rect 1301 5538 1367 5541
rect 0 5536 1367 5538
rect 0 5480 1306 5536
rect 1362 5480 1367 5536
rect 0 5478 1367 5480
rect 0 5448 800 5478
rect 1301 5475 1367 5478
rect 10593 5538 10659 5541
rect 11198 5538 11998 5568
rect 10593 5536 11998 5538
rect 10593 5480 10598 5536
rect 10654 5480 11998 5536
rect 10593 5478 11998 5480
rect 10593 5475 10659 5478
rect 2825 5472 3141 5473
rect 2825 5408 2831 5472
rect 2895 5408 2911 5472
rect 2975 5408 2991 5472
rect 3055 5408 3071 5472
rect 3135 5408 3141 5472
rect 2825 5407 3141 5408
rect 5263 5472 5579 5473
rect 5263 5408 5269 5472
rect 5333 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5579 5472
rect 5263 5407 5579 5408
rect 7701 5472 8017 5473
rect 7701 5408 7707 5472
rect 7771 5408 7787 5472
rect 7851 5408 7867 5472
rect 7931 5408 7947 5472
rect 8011 5408 8017 5472
rect 7701 5407 8017 5408
rect 10139 5472 10455 5473
rect 10139 5408 10145 5472
rect 10209 5408 10225 5472
rect 10289 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10455 5472
rect 11198 5448 11998 5478
rect 10139 5407 10455 5408
rect 6821 5266 6887 5269
rect 7465 5266 7531 5269
rect 6821 5264 7531 5266
rect 6821 5208 6826 5264
rect 6882 5208 7470 5264
rect 7526 5208 7531 5264
rect 6821 5206 7531 5208
rect 6821 5203 6887 5206
rect 7465 5203 7531 5206
rect 2165 4928 2481 4929
rect 0 4858 800 4888
rect 2165 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2481 4928
rect 2165 4863 2481 4864
rect 4603 4928 4919 4929
rect 4603 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4919 4928
rect 4603 4863 4919 4864
rect 7041 4928 7357 4929
rect 7041 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7357 4928
rect 7041 4863 7357 4864
rect 9479 4928 9795 4929
rect 9479 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9795 4928
rect 9479 4863 9795 4864
rect 10501 4858 10567 4861
rect 11198 4858 11998 4888
rect 0 4768 858 4858
rect 10501 4856 11998 4858
rect 10501 4800 10506 4856
rect 10562 4800 11998 4856
rect 10501 4798 11998 4800
rect 10501 4795 10567 4798
rect 11198 4768 11998 4798
rect 798 4725 858 4768
rect 798 4720 907 4725
rect 798 4664 846 4720
rect 902 4664 907 4720
rect 798 4662 907 4664
rect 841 4659 907 4662
rect 2825 4384 3141 4385
rect 2825 4320 2831 4384
rect 2895 4320 2911 4384
rect 2975 4320 2991 4384
rect 3055 4320 3071 4384
rect 3135 4320 3141 4384
rect 2825 4319 3141 4320
rect 5263 4384 5579 4385
rect 5263 4320 5269 4384
rect 5333 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5579 4384
rect 5263 4319 5579 4320
rect 7701 4384 8017 4385
rect 7701 4320 7707 4384
rect 7771 4320 7787 4384
rect 7851 4320 7867 4384
rect 7931 4320 7947 4384
rect 8011 4320 8017 4384
rect 7701 4319 8017 4320
rect 10139 4384 10455 4385
rect 10139 4320 10145 4384
rect 10209 4320 10225 4384
rect 10289 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10455 4384
rect 10139 4319 10455 4320
rect 2165 3840 2481 3841
rect 2165 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2481 3840
rect 2165 3775 2481 3776
rect 4603 3840 4919 3841
rect 4603 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4919 3840
rect 4603 3775 4919 3776
rect 7041 3840 7357 3841
rect 7041 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7357 3840
rect 7041 3775 7357 3776
rect 9479 3840 9795 3841
rect 9479 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9795 3840
rect 9479 3775 9795 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 2589 3634 2655 3637
rect 3509 3634 3575 3637
rect 7465 3634 7531 3637
rect 2589 3632 7531 3634
rect 2589 3576 2594 3632
rect 2650 3576 3514 3632
rect 3570 3576 7470 3632
rect 7526 3576 7531 3632
rect 2589 3574 7531 3576
rect 2589 3571 2655 3574
rect 3509 3571 3575 3574
rect 7465 3571 7531 3574
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 0 3408 800 3438
rect 2825 3296 3141 3297
rect 2825 3232 2831 3296
rect 2895 3232 2911 3296
rect 2975 3232 2991 3296
rect 3055 3232 3071 3296
rect 3135 3232 3141 3296
rect 2825 3231 3141 3232
rect 5263 3296 5579 3297
rect 5263 3232 5269 3296
rect 5333 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5579 3296
rect 5263 3231 5579 3232
rect 7701 3296 8017 3297
rect 7701 3232 7707 3296
rect 7771 3232 7787 3296
rect 7851 3232 7867 3296
rect 7931 3232 7947 3296
rect 8011 3232 8017 3296
rect 7701 3231 8017 3232
rect 10139 3296 10455 3297
rect 10139 3232 10145 3296
rect 10209 3232 10225 3296
rect 10289 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10455 3296
rect 10139 3231 10455 3232
rect 4061 3090 4127 3093
rect 7097 3090 7163 3093
rect 4061 3088 7163 3090
rect 4061 3032 4066 3088
rect 4122 3032 7102 3088
rect 7158 3032 7163 3088
rect 4061 3030 7163 3032
rect 4061 3027 4127 3030
rect 7097 3027 7163 3030
rect 2165 2752 2481 2753
rect 2165 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2481 2752
rect 2165 2687 2481 2688
rect 4603 2752 4919 2753
rect 4603 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4919 2752
rect 4603 2687 4919 2688
rect 7041 2752 7357 2753
rect 7041 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7357 2752
rect 7041 2687 7357 2688
rect 9479 2752 9795 2753
rect 9479 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9795 2752
rect 9479 2687 9795 2688
rect 2825 2208 3141 2209
rect 2825 2144 2831 2208
rect 2895 2144 2911 2208
rect 2975 2144 2991 2208
rect 3055 2144 3071 2208
rect 3135 2144 3141 2208
rect 2825 2143 3141 2144
rect 5263 2208 5579 2209
rect 5263 2144 5269 2208
rect 5333 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5579 2208
rect 5263 2143 5579 2144
rect 7701 2208 8017 2209
rect 7701 2144 7707 2208
rect 7771 2144 7787 2208
rect 7851 2144 7867 2208
rect 7931 2144 7947 2208
rect 8011 2144 8017 2208
rect 7701 2143 8017 2144
rect 10139 2208 10455 2209
rect 10139 2144 10145 2208
rect 10209 2144 10225 2208
rect 10289 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10455 2208
rect 10139 2143 10455 2144
<< via3 >>
rect 2171 11452 2235 11456
rect 2171 11396 2175 11452
rect 2175 11396 2231 11452
rect 2231 11396 2235 11452
rect 2171 11392 2235 11396
rect 2251 11452 2315 11456
rect 2251 11396 2255 11452
rect 2255 11396 2311 11452
rect 2311 11396 2315 11452
rect 2251 11392 2315 11396
rect 2331 11452 2395 11456
rect 2331 11396 2335 11452
rect 2335 11396 2391 11452
rect 2391 11396 2395 11452
rect 2331 11392 2395 11396
rect 2411 11452 2475 11456
rect 2411 11396 2415 11452
rect 2415 11396 2471 11452
rect 2471 11396 2475 11452
rect 2411 11392 2475 11396
rect 4609 11452 4673 11456
rect 4609 11396 4613 11452
rect 4613 11396 4669 11452
rect 4669 11396 4673 11452
rect 4609 11392 4673 11396
rect 4689 11452 4753 11456
rect 4689 11396 4693 11452
rect 4693 11396 4749 11452
rect 4749 11396 4753 11452
rect 4689 11392 4753 11396
rect 4769 11452 4833 11456
rect 4769 11396 4773 11452
rect 4773 11396 4829 11452
rect 4829 11396 4833 11452
rect 4769 11392 4833 11396
rect 4849 11452 4913 11456
rect 4849 11396 4853 11452
rect 4853 11396 4909 11452
rect 4909 11396 4913 11452
rect 4849 11392 4913 11396
rect 7047 11452 7111 11456
rect 7047 11396 7051 11452
rect 7051 11396 7107 11452
rect 7107 11396 7111 11452
rect 7047 11392 7111 11396
rect 7127 11452 7191 11456
rect 7127 11396 7131 11452
rect 7131 11396 7187 11452
rect 7187 11396 7191 11452
rect 7127 11392 7191 11396
rect 7207 11452 7271 11456
rect 7207 11396 7211 11452
rect 7211 11396 7267 11452
rect 7267 11396 7271 11452
rect 7207 11392 7271 11396
rect 7287 11452 7351 11456
rect 7287 11396 7291 11452
rect 7291 11396 7347 11452
rect 7347 11396 7351 11452
rect 7287 11392 7351 11396
rect 9485 11452 9549 11456
rect 9485 11396 9489 11452
rect 9489 11396 9545 11452
rect 9545 11396 9549 11452
rect 9485 11392 9549 11396
rect 9565 11452 9629 11456
rect 9565 11396 9569 11452
rect 9569 11396 9625 11452
rect 9625 11396 9629 11452
rect 9565 11392 9629 11396
rect 9645 11452 9709 11456
rect 9645 11396 9649 11452
rect 9649 11396 9705 11452
rect 9705 11396 9709 11452
rect 9645 11392 9709 11396
rect 9725 11452 9789 11456
rect 9725 11396 9729 11452
rect 9729 11396 9785 11452
rect 9785 11396 9789 11452
rect 9725 11392 9789 11396
rect 2831 10908 2895 10912
rect 2831 10852 2835 10908
rect 2835 10852 2891 10908
rect 2891 10852 2895 10908
rect 2831 10848 2895 10852
rect 2911 10908 2975 10912
rect 2911 10852 2915 10908
rect 2915 10852 2971 10908
rect 2971 10852 2975 10908
rect 2911 10848 2975 10852
rect 2991 10908 3055 10912
rect 2991 10852 2995 10908
rect 2995 10852 3051 10908
rect 3051 10852 3055 10908
rect 2991 10848 3055 10852
rect 3071 10908 3135 10912
rect 3071 10852 3075 10908
rect 3075 10852 3131 10908
rect 3131 10852 3135 10908
rect 3071 10848 3135 10852
rect 5269 10908 5333 10912
rect 5269 10852 5273 10908
rect 5273 10852 5329 10908
rect 5329 10852 5333 10908
rect 5269 10848 5333 10852
rect 5349 10908 5413 10912
rect 5349 10852 5353 10908
rect 5353 10852 5409 10908
rect 5409 10852 5413 10908
rect 5349 10848 5413 10852
rect 5429 10908 5493 10912
rect 5429 10852 5433 10908
rect 5433 10852 5489 10908
rect 5489 10852 5493 10908
rect 5429 10848 5493 10852
rect 5509 10908 5573 10912
rect 5509 10852 5513 10908
rect 5513 10852 5569 10908
rect 5569 10852 5573 10908
rect 5509 10848 5573 10852
rect 7707 10908 7771 10912
rect 7707 10852 7711 10908
rect 7711 10852 7767 10908
rect 7767 10852 7771 10908
rect 7707 10848 7771 10852
rect 7787 10908 7851 10912
rect 7787 10852 7791 10908
rect 7791 10852 7847 10908
rect 7847 10852 7851 10908
rect 7787 10848 7851 10852
rect 7867 10908 7931 10912
rect 7867 10852 7871 10908
rect 7871 10852 7927 10908
rect 7927 10852 7931 10908
rect 7867 10848 7931 10852
rect 7947 10908 8011 10912
rect 7947 10852 7951 10908
rect 7951 10852 8007 10908
rect 8007 10852 8011 10908
rect 7947 10848 8011 10852
rect 10145 10908 10209 10912
rect 10145 10852 10149 10908
rect 10149 10852 10205 10908
rect 10205 10852 10209 10908
rect 10145 10848 10209 10852
rect 10225 10908 10289 10912
rect 10225 10852 10229 10908
rect 10229 10852 10285 10908
rect 10285 10852 10289 10908
rect 10225 10848 10289 10852
rect 10305 10908 10369 10912
rect 10305 10852 10309 10908
rect 10309 10852 10365 10908
rect 10365 10852 10369 10908
rect 10305 10848 10369 10852
rect 10385 10908 10449 10912
rect 10385 10852 10389 10908
rect 10389 10852 10445 10908
rect 10445 10852 10449 10908
rect 10385 10848 10449 10852
rect 2171 10364 2235 10368
rect 2171 10308 2175 10364
rect 2175 10308 2231 10364
rect 2231 10308 2235 10364
rect 2171 10304 2235 10308
rect 2251 10364 2315 10368
rect 2251 10308 2255 10364
rect 2255 10308 2311 10364
rect 2311 10308 2315 10364
rect 2251 10304 2315 10308
rect 2331 10364 2395 10368
rect 2331 10308 2335 10364
rect 2335 10308 2391 10364
rect 2391 10308 2395 10364
rect 2331 10304 2395 10308
rect 2411 10364 2475 10368
rect 2411 10308 2415 10364
rect 2415 10308 2471 10364
rect 2471 10308 2475 10364
rect 2411 10304 2475 10308
rect 4609 10364 4673 10368
rect 4609 10308 4613 10364
rect 4613 10308 4669 10364
rect 4669 10308 4673 10364
rect 4609 10304 4673 10308
rect 4689 10364 4753 10368
rect 4689 10308 4693 10364
rect 4693 10308 4749 10364
rect 4749 10308 4753 10364
rect 4689 10304 4753 10308
rect 4769 10364 4833 10368
rect 4769 10308 4773 10364
rect 4773 10308 4829 10364
rect 4829 10308 4833 10364
rect 4769 10304 4833 10308
rect 4849 10364 4913 10368
rect 4849 10308 4853 10364
rect 4853 10308 4909 10364
rect 4909 10308 4913 10364
rect 4849 10304 4913 10308
rect 7047 10364 7111 10368
rect 7047 10308 7051 10364
rect 7051 10308 7107 10364
rect 7107 10308 7111 10364
rect 7047 10304 7111 10308
rect 7127 10364 7191 10368
rect 7127 10308 7131 10364
rect 7131 10308 7187 10364
rect 7187 10308 7191 10364
rect 7127 10304 7191 10308
rect 7207 10364 7271 10368
rect 7207 10308 7211 10364
rect 7211 10308 7267 10364
rect 7267 10308 7271 10364
rect 7207 10304 7271 10308
rect 7287 10364 7351 10368
rect 7287 10308 7291 10364
rect 7291 10308 7347 10364
rect 7347 10308 7351 10364
rect 7287 10304 7351 10308
rect 9485 10364 9549 10368
rect 9485 10308 9489 10364
rect 9489 10308 9545 10364
rect 9545 10308 9549 10364
rect 9485 10304 9549 10308
rect 9565 10364 9629 10368
rect 9565 10308 9569 10364
rect 9569 10308 9625 10364
rect 9625 10308 9629 10364
rect 9565 10304 9629 10308
rect 9645 10364 9709 10368
rect 9645 10308 9649 10364
rect 9649 10308 9705 10364
rect 9705 10308 9709 10364
rect 9645 10304 9709 10308
rect 9725 10364 9789 10368
rect 9725 10308 9729 10364
rect 9729 10308 9785 10364
rect 9785 10308 9789 10364
rect 9725 10304 9789 10308
rect 2831 9820 2895 9824
rect 2831 9764 2835 9820
rect 2835 9764 2891 9820
rect 2891 9764 2895 9820
rect 2831 9760 2895 9764
rect 2911 9820 2975 9824
rect 2911 9764 2915 9820
rect 2915 9764 2971 9820
rect 2971 9764 2975 9820
rect 2911 9760 2975 9764
rect 2991 9820 3055 9824
rect 2991 9764 2995 9820
rect 2995 9764 3051 9820
rect 3051 9764 3055 9820
rect 2991 9760 3055 9764
rect 3071 9820 3135 9824
rect 3071 9764 3075 9820
rect 3075 9764 3131 9820
rect 3131 9764 3135 9820
rect 3071 9760 3135 9764
rect 5269 9820 5333 9824
rect 5269 9764 5273 9820
rect 5273 9764 5329 9820
rect 5329 9764 5333 9820
rect 5269 9760 5333 9764
rect 5349 9820 5413 9824
rect 5349 9764 5353 9820
rect 5353 9764 5409 9820
rect 5409 9764 5413 9820
rect 5349 9760 5413 9764
rect 5429 9820 5493 9824
rect 5429 9764 5433 9820
rect 5433 9764 5489 9820
rect 5489 9764 5493 9820
rect 5429 9760 5493 9764
rect 5509 9820 5573 9824
rect 5509 9764 5513 9820
rect 5513 9764 5569 9820
rect 5569 9764 5573 9820
rect 5509 9760 5573 9764
rect 7707 9820 7771 9824
rect 7707 9764 7711 9820
rect 7711 9764 7767 9820
rect 7767 9764 7771 9820
rect 7707 9760 7771 9764
rect 7787 9820 7851 9824
rect 7787 9764 7791 9820
rect 7791 9764 7847 9820
rect 7847 9764 7851 9820
rect 7787 9760 7851 9764
rect 7867 9820 7931 9824
rect 7867 9764 7871 9820
rect 7871 9764 7927 9820
rect 7927 9764 7931 9820
rect 7867 9760 7931 9764
rect 7947 9820 8011 9824
rect 7947 9764 7951 9820
rect 7951 9764 8007 9820
rect 8007 9764 8011 9820
rect 7947 9760 8011 9764
rect 10145 9820 10209 9824
rect 10145 9764 10149 9820
rect 10149 9764 10205 9820
rect 10205 9764 10209 9820
rect 10145 9760 10209 9764
rect 10225 9820 10289 9824
rect 10225 9764 10229 9820
rect 10229 9764 10285 9820
rect 10285 9764 10289 9820
rect 10225 9760 10289 9764
rect 10305 9820 10369 9824
rect 10305 9764 10309 9820
rect 10309 9764 10365 9820
rect 10365 9764 10369 9820
rect 10305 9760 10369 9764
rect 10385 9820 10449 9824
rect 10385 9764 10389 9820
rect 10389 9764 10445 9820
rect 10445 9764 10449 9820
rect 10385 9760 10449 9764
rect 2171 9276 2235 9280
rect 2171 9220 2175 9276
rect 2175 9220 2231 9276
rect 2231 9220 2235 9276
rect 2171 9216 2235 9220
rect 2251 9276 2315 9280
rect 2251 9220 2255 9276
rect 2255 9220 2311 9276
rect 2311 9220 2315 9276
rect 2251 9216 2315 9220
rect 2331 9276 2395 9280
rect 2331 9220 2335 9276
rect 2335 9220 2391 9276
rect 2391 9220 2395 9276
rect 2331 9216 2395 9220
rect 2411 9276 2475 9280
rect 2411 9220 2415 9276
rect 2415 9220 2471 9276
rect 2471 9220 2475 9276
rect 2411 9216 2475 9220
rect 4609 9276 4673 9280
rect 4609 9220 4613 9276
rect 4613 9220 4669 9276
rect 4669 9220 4673 9276
rect 4609 9216 4673 9220
rect 4689 9276 4753 9280
rect 4689 9220 4693 9276
rect 4693 9220 4749 9276
rect 4749 9220 4753 9276
rect 4689 9216 4753 9220
rect 4769 9276 4833 9280
rect 4769 9220 4773 9276
rect 4773 9220 4829 9276
rect 4829 9220 4833 9276
rect 4769 9216 4833 9220
rect 4849 9276 4913 9280
rect 4849 9220 4853 9276
rect 4853 9220 4909 9276
rect 4909 9220 4913 9276
rect 4849 9216 4913 9220
rect 7047 9276 7111 9280
rect 7047 9220 7051 9276
rect 7051 9220 7107 9276
rect 7107 9220 7111 9276
rect 7047 9216 7111 9220
rect 7127 9276 7191 9280
rect 7127 9220 7131 9276
rect 7131 9220 7187 9276
rect 7187 9220 7191 9276
rect 7127 9216 7191 9220
rect 7207 9276 7271 9280
rect 7207 9220 7211 9276
rect 7211 9220 7267 9276
rect 7267 9220 7271 9276
rect 7207 9216 7271 9220
rect 7287 9276 7351 9280
rect 7287 9220 7291 9276
rect 7291 9220 7347 9276
rect 7347 9220 7351 9276
rect 7287 9216 7351 9220
rect 9485 9276 9549 9280
rect 9485 9220 9489 9276
rect 9489 9220 9545 9276
rect 9545 9220 9549 9276
rect 9485 9216 9549 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 2831 8732 2895 8736
rect 2831 8676 2835 8732
rect 2835 8676 2891 8732
rect 2891 8676 2895 8732
rect 2831 8672 2895 8676
rect 2911 8732 2975 8736
rect 2911 8676 2915 8732
rect 2915 8676 2971 8732
rect 2971 8676 2975 8732
rect 2911 8672 2975 8676
rect 2991 8732 3055 8736
rect 2991 8676 2995 8732
rect 2995 8676 3051 8732
rect 3051 8676 3055 8732
rect 2991 8672 3055 8676
rect 3071 8732 3135 8736
rect 3071 8676 3075 8732
rect 3075 8676 3131 8732
rect 3131 8676 3135 8732
rect 3071 8672 3135 8676
rect 5269 8732 5333 8736
rect 5269 8676 5273 8732
rect 5273 8676 5329 8732
rect 5329 8676 5333 8732
rect 5269 8672 5333 8676
rect 5349 8732 5413 8736
rect 5349 8676 5353 8732
rect 5353 8676 5409 8732
rect 5409 8676 5413 8732
rect 5349 8672 5413 8676
rect 5429 8732 5493 8736
rect 5429 8676 5433 8732
rect 5433 8676 5489 8732
rect 5489 8676 5493 8732
rect 5429 8672 5493 8676
rect 5509 8732 5573 8736
rect 5509 8676 5513 8732
rect 5513 8676 5569 8732
rect 5569 8676 5573 8732
rect 5509 8672 5573 8676
rect 7707 8732 7771 8736
rect 7707 8676 7711 8732
rect 7711 8676 7767 8732
rect 7767 8676 7771 8732
rect 7707 8672 7771 8676
rect 7787 8732 7851 8736
rect 7787 8676 7791 8732
rect 7791 8676 7847 8732
rect 7847 8676 7851 8732
rect 7787 8672 7851 8676
rect 7867 8732 7931 8736
rect 7867 8676 7871 8732
rect 7871 8676 7927 8732
rect 7927 8676 7931 8732
rect 7867 8672 7931 8676
rect 7947 8732 8011 8736
rect 7947 8676 7951 8732
rect 7951 8676 8007 8732
rect 8007 8676 8011 8732
rect 7947 8672 8011 8676
rect 10145 8732 10209 8736
rect 10145 8676 10149 8732
rect 10149 8676 10205 8732
rect 10205 8676 10209 8732
rect 10145 8672 10209 8676
rect 10225 8732 10289 8736
rect 10225 8676 10229 8732
rect 10229 8676 10285 8732
rect 10285 8676 10289 8732
rect 10225 8672 10289 8676
rect 10305 8732 10369 8736
rect 10305 8676 10309 8732
rect 10309 8676 10365 8732
rect 10365 8676 10369 8732
rect 10305 8672 10369 8676
rect 10385 8732 10449 8736
rect 10385 8676 10389 8732
rect 10389 8676 10445 8732
rect 10445 8676 10449 8732
rect 10385 8672 10449 8676
rect 2171 8188 2235 8192
rect 2171 8132 2175 8188
rect 2175 8132 2231 8188
rect 2231 8132 2235 8188
rect 2171 8128 2235 8132
rect 2251 8188 2315 8192
rect 2251 8132 2255 8188
rect 2255 8132 2311 8188
rect 2311 8132 2315 8188
rect 2251 8128 2315 8132
rect 2331 8188 2395 8192
rect 2331 8132 2335 8188
rect 2335 8132 2391 8188
rect 2391 8132 2395 8188
rect 2331 8128 2395 8132
rect 2411 8188 2475 8192
rect 2411 8132 2415 8188
rect 2415 8132 2471 8188
rect 2471 8132 2475 8188
rect 2411 8128 2475 8132
rect 4609 8188 4673 8192
rect 4609 8132 4613 8188
rect 4613 8132 4669 8188
rect 4669 8132 4673 8188
rect 4609 8128 4673 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 7047 8188 7111 8192
rect 7047 8132 7051 8188
rect 7051 8132 7107 8188
rect 7107 8132 7111 8188
rect 7047 8128 7111 8132
rect 7127 8188 7191 8192
rect 7127 8132 7131 8188
rect 7131 8132 7187 8188
rect 7187 8132 7191 8188
rect 7127 8128 7191 8132
rect 7207 8188 7271 8192
rect 7207 8132 7211 8188
rect 7211 8132 7267 8188
rect 7267 8132 7271 8188
rect 7207 8128 7271 8132
rect 7287 8188 7351 8192
rect 7287 8132 7291 8188
rect 7291 8132 7347 8188
rect 7347 8132 7351 8188
rect 7287 8128 7351 8132
rect 9485 8188 9549 8192
rect 9485 8132 9489 8188
rect 9489 8132 9545 8188
rect 9545 8132 9549 8188
rect 9485 8128 9549 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 2831 7644 2895 7648
rect 2831 7588 2835 7644
rect 2835 7588 2891 7644
rect 2891 7588 2895 7644
rect 2831 7584 2895 7588
rect 2911 7644 2975 7648
rect 2911 7588 2915 7644
rect 2915 7588 2971 7644
rect 2971 7588 2975 7644
rect 2911 7584 2975 7588
rect 2991 7644 3055 7648
rect 2991 7588 2995 7644
rect 2995 7588 3051 7644
rect 3051 7588 3055 7644
rect 2991 7584 3055 7588
rect 3071 7644 3135 7648
rect 3071 7588 3075 7644
rect 3075 7588 3131 7644
rect 3131 7588 3135 7644
rect 3071 7584 3135 7588
rect 5269 7644 5333 7648
rect 5269 7588 5273 7644
rect 5273 7588 5329 7644
rect 5329 7588 5333 7644
rect 5269 7584 5333 7588
rect 5349 7644 5413 7648
rect 5349 7588 5353 7644
rect 5353 7588 5409 7644
rect 5409 7588 5413 7644
rect 5349 7584 5413 7588
rect 5429 7644 5493 7648
rect 5429 7588 5433 7644
rect 5433 7588 5489 7644
rect 5489 7588 5493 7644
rect 5429 7584 5493 7588
rect 5509 7644 5573 7648
rect 5509 7588 5513 7644
rect 5513 7588 5569 7644
rect 5569 7588 5573 7644
rect 5509 7584 5573 7588
rect 7707 7644 7771 7648
rect 7707 7588 7711 7644
rect 7711 7588 7767 7644
rect 7767 7588 7771 7644
rect 7707 7584 7771 7588
rect 7787 7644 7851 7648
rect 7787 7588 7791 7644
rect 7791 7588 7847 7644
rect 7847 7588 7851 7644
rect 7787 7584 7851 7588
rect 7867 7644 7931 7648
rect 7867 7588 7871 7644
rect 7871 7588 7927 7644
rect 7927 7588 7931 7644
rect 7867 7584 7931 7588
rect 7947 7644 8011 7648
rect 7947 7588 7951 7644
rect 7951 7588 8007 7644
rect 8007 7588 8011 7644
rect 7947 7584 8011 7588
rect 10145 7644 10209 7648
rect 10145 7588 10149 7644
rect 10149 7588 10205 7644
rect 10205 7588 10209 7644
rect 10145 7584 10209 7588
rect 10225 7644 10289 7648
rect 10225 7588 10229 7644
rect 10229 7588 10285 7644
rect 10285 7588 10289 7644
rect 10225 7584 10289 7588
rect 10305 7644 10369 7648
rect 10305 7588 10309 7644
rect 10309 7588 10365 7644
rect 10365 7588 10369 7644
rect 10305 7584 10369 7588
rect 10385 7644 10449 7648
rect 10385 7588 10389 7644
rect 10389 7588 10445 7644
rect 10445 7588 10449 7644
rect 10385 7584 10449 7588
rect 2171 7100 2235 7104
rect 2171 7044 2175 7100
rect 2175 7044 2231 7100
rect 2231 7044 2235 7100
rect 2171 7040 2235 7044
rect 2251 7100 2315 7104
rect 2251 7044 2255 7100
rect 2255 7044 2311 7100
rect 2311 7044 2315 7100
rect 2251 7040 2315 7044
rect 2331 7100 2395 7104
rect 2331 7044 2335 7100
rect 2335 7044 2391 7100
rect 2391 7044 2395 7100
rect 2331 7040 2395 7044
rect 2411 7100 2475 7104
rect 2411 7044 2415 7100
rect 2415 7044 2471 7100
rect 2471 7044 2475 7100
rect 2411 7040 2475 7044
rect 4609 7100 4673 7104
rect 4609 7044 4613 7100
rect 4613 7044 4669 7100
rect 4669 7044 4673 7100
rect 4609 7040 4673 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 7047 7100 7111 7104
rect 7047 7044 7051 7100
rect 7051 7044 7107 7100
rect 7107 7044 7111 7100
rect 7047 7040 7111 7044
rect 7127 7100 7191 7104
rect 7127 7044 7131 7100
rect 7131 7044 7187 7100
rect 7187 7044 7191 7100
rect 7127 7040 7191 7044
rect 7207 7100 7271 7104
rect 7207 7044 7211 7100
rect 7211 7044 7267 7100
rect 7267 7044 7271 7100
rect 7207 7040 7271 7044
rect 7287 7100 7351 7104
rect 7287 7044 7291 7100
rect 7291 7044 7347 7100
rect 7347 7044 7351 7100
rect 7287 7040 7351 7044
rect 9485 7100 9549 7104
rect 9485 7044 9489 7100
rect 9489 7044 9545 7100
rect 9545 7044 9549 7100
rect 9485 7040 9549 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 2831 6556 2895 6560
rect 2831 6500 2835 6556
rect 2835 6500 2891 6556
rect 2891 6500 2895 6556
rect 2831 6496 2895 6500
rect 2911 6556 2975 6560
rect 2911 6500 2915 6556
rect 2915 6500 2971 6556
rect 2971 6500 2975 6556
rect 2911 6496 2975 6500
rect 2991 6556 3055 6560
rect 2991 6500 2995 6556
rect 2995 6500 3051 6556
rect 3051 6500 3055 6556
rect 2991 6496 3055 6500
rect 3071 6556 3135 6560
rect 3071 6500 3075 6556
rect 3075 6500 3131 6556
rect 3131 6500 3135 6556
rect 3071 6496 3135 6500
rect 5269 6556 5333 6560
rect 5269 6500 5273 6556
rect 5273 6500 5329 6556
rect 5329 6500 5333 6556
rect 5269 6496 5333 6500
rect 5349 6556 5413 6560
rect 5349 6500 5353 6556
rect 5353 6500 5409 6556
rect 5409 6500 5413 6556
rect 5349 6496 5413 6500
rect 5429 6556 5493 6560
rect 5429 6500 5433 6556
rect 5433 6500 5489 6556
rect 5489 6500 5493 6556
rect 5429 6496 5493 6500
rect 5509 6556 5573 6560
rect 5509 6500 5513 6556
rect 5513 6500 5569 6556
rect 5569 6500 5573 6556
rect 5509 6496 5573 6500
rect 7707 6556 7771 6560
rect 7707 6500 7711 6556
rect 7711 6500 7767 6556
rect 7767 6500 7771 6556
rect 7707 6496 7771 6500
rect 7787 6556 7851 6560
rect 7787 6500 7791 6556
rect 7791 6500 7847 6556
rect 7847 6500 7851 6556
rect 7787 6496 7851 6500
rect 7867 6556 7931 6560
rect 7867 6500 7871 6556
rect 7871 6500 7927 6556
rect 7927 6500 7931 6556
rect 7867 6496 7931 6500
rect 7947 6556 8011 6560
rect 7947 6500 7951 6556
rect 7951 6500 8007 6556
rect 8007 6500 8011 6556
rect 7947 6496 8011 6500
rect 10145 6556 10209 6560
rect 10145 6500 10149 6556
rect 10149 6500 10205 6556
rect 10205 6500 10209 6556
rect 10145 6496 10209 6500
rect 10225 6556 10289 6560
rect 10225 6500 10229 6556
rect 10229 6500 10285 6556
rect 10285 6500 10289 6556
rect 10225 6496 10289 6500
rect 10305 6556 10369 6560
rect 10305 6500 10309 6556
rect 10309 6500 10365 6556
rect 10365 6500 10369 6556
rect 10305 6496 10369 6500
rect 10385 6556 10449 6560
rect 10385 6500 10389 6556
rect 10389 6500 10445 6556
rect 10445 6500 10449 6556
rect 10385 6496 10449 6500
rect 2171 6012 2235 6016
rect 2171 5956 2175 6012
rect 2175 5956 2231 6012
rect 2231 5956 2235 6012
rect 2171 5952 2235 5956
rect 2251 6012 2315 6016
rect 2251 5956 2255 6012
rect 2255 5956 2311 6012
rect 2311 5956 2315 6012
rect 2251 5952 2315 5956
rect 2331 6012 2395 6016
rect 2331 5956 2335 6012
rect 2335 5956 2391 6012
rect 2391 5956 2395 6012
rect 2331 5952 2395 5956
rect 2411 6012 2475 6016
rect 2411 5956 2415 6012
rect 2415 5956 2471 6012
rect 2471 5956 2475 6012
rect 2411 5952 2475 5956
rect 4609 6012 4673 6016
rect 4609 5956 4613 6012
rect 4613 5956 4669 6012
rect 4669 5956 4673 6012
rect 4609 5952 4673 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 7047 6012 7111 6016
rect 7047 5956 7051 6012
rect 7051 5956 7107 6012
rect 7107 5956 7111 6012
rect 7047 5952 7111 5956
rect 7127 6012 7191 6016
rect 7127 5956 7131 6012
rect 7131 5956 7187 6012
rect 7187 5956 7191 6012
rect 7127 5952 7191 5956
rect 7207 6012 7271 6016
rect 7207 5956 7211 6012
rect 7211 5956 7267 6012
rect 7267 5956 7271 6012
rect 7207 5952 7271 5956
rect 7287 6012 7351 6016
rect 7287 5956 7291 6012
rect 7291 5956 7347 6012
rect 7347 5956 7351 6012
rect 7287 5952 7351 5956
rect 9485 6012 9549 6016
rect 9485 5956 9489 6012
rect 9489 5956 9545 6012
rect 9545 5956 9549 6012
rect 9485 5952 9549 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 2831 5468 2895 5472
rect 2831 5412 2835 5468
rect 2835 5412 2891 5468
rect 2891 5412 2895 5468
rect 2831 5408 2895 5412
rect 2911 5468 2975 5472
rect 2911 5412 2915 5468
rect 2915 5412 2971 5468
rect 2971 5412 2975 5468
rect 2911 5408 2975 5412
rect 2991 5468 3055 5472
rect 2991 5412 2995 5468
rect 2995 5412 3051 5468
rect 3051 5412 3055 5468
rect 2991 5408 3055 5412
rect 3071 5468 3135 5472
rect 3071 5412 3075 5468
rect 3075 5412 3131 5468
rect 3131 5412 3135 5468
rect 3071 5408 3135 5412
rect 5269 5468 5333 5472
rect 5269 5412 5273 5468
rect 5273 5412 5329 5468
rect 5329 5412 5333 5468
rect 5269 5408 5333 5412
rect 5349 5468 5413 5472
rect 5349 5412 5353 5468
rect 5353 5412 5409 5468
rect 5409 5412 5413 5468
rect 5349 5408 5413 5412
rect 5429 5468 5493 5472
rect 5429 5412 5433 5468
rect 5433 5412 5489 5468
rect 5489 5412 5493 5468
rect 5429 5408 5493 5412
rect 5509 5468 5573 5472
rect 5509 5412 5513 5468
rect 5513 5412 5569 5468
rect 5569 5412 5573 5468
rect 5509 5408 5573 5412
rect 7707 5468 7771 5472
rect 7707 5412 7711 5468
rect 7711 5412 7767 5468
rect 7767 5412 7771 5468
rect 7707 5408 7771 5412
rect 7787 5468 7851 5472
rect 7787 5412 7791 5468
rect 7791 5412 7847 5468
rect 7847 5412 7851 5468
rect 7787 5408 7851 5412
rect 7867 5468 7931 5472
rect 7867 5412 7871 5468
rect 7871 5412 7927 5468
rect 7927 5412 7931 5468
rect 7867 5408 7931 5412
rect 7947 5468 8011 5472
rect 7947 5412 7951 5468
rect 7951 5412 8007 5468
rect 8007 5412 8011 5468
rect 7947 5408 8011 5412
rect 10145 5468 10209 5472
rect 10145 5412 10149 5468
rect 10149 5412 10205 5468
rect 10205 5412 10209 5468
rect 10145 5408 10209 5412
rect 10225 5468 10289 5472
rect 10225 5412 10229 5468
rect 10229 5412 10285 5468
rect 10285 5412 10289 5468
rect 10225 5408 10289 5412
rect 10305 5468 10369 5472
rect 10305 5412 10309 5468
rect 10309 5412 10365 5468
rect 10365 5412 10369 5468
rect 10305 5408 10369 5412
rect 10385 5468 10449 5472
rect 10385 5412 10389 5468
rect 10389 5412 10445 5468
rect 10445 5412 10449 5468
rect 10385 5408 10449 5412
rect 2171 4924 2235 4928
rect 2171 4868 2175 4924
rect 2175 4868 2231 4924
rect 2231 4868 2235 4924
rect 2171 4864 2235 4868
rect 2251 4924 2315 4928
rect 2251 4868 2255 4924
rect 2255 4868 2311 4924
rect 2311 4868 2315 4924
rect 2251 4864 2315 4868
rect 2331 4924 2395 4928
rect 2331 4868 2335 4924
rect 2335 4868 2391 4924
rect 2391 4868 2395 4924
rect 2331 4864 2395 4868
rect 2411 4924 2475 4928
rect 2411 4868 2415 4924
rect 2415 4868 2471 4924
rect 2471 4868 2475 4924
rect 2411 4864 2475 4868
rect 4609 4924 4673 4928
rect 4609 4868 4613 4924
rect 4613 4868 4669 4924
rect 4669 4868 4673 4924
rect 4609 4864 4673 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 7047 4924 7111 4928
rect 7047 4868 7051 4924
rect 7051 4868 7107 4924
rect 7107 4868 7111 4924
rect 7047 4864 7111 4868
rect 7127 4924 7191 4928
rect 7127 4868 7131 4924
rect 7131 4868 7187 4924
rect 7187 4868 7191 4924
rect 7127 4864 7191 4868
rect 7207 4924 7271 4928
rect 7207 4868 7211 4924
rect 7211 4868 7267 4924
rect 7267 4868 7271 4924
rect 7207 4864 7271 4868
rect 7287 4924 7351 4928
rect 7287 4868 7291 4924
rect 7291 4868 7347 4924
rect 7347 4868 7351 4924
rect 7287 4864 7351 4868
rect 9485 4924 9549 4928
rect 9485 4868 9489 4924
rect 9489 4868 9545 4924
rect 9545 4868 9549 4924
rect 9485 4864 9549 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 2831 4380 2895 4384
rect 2831 4324 2835 4380
rect 2835 4324 2891 4380
rect 2891 4324 2895 4380
rect 2831 4320 2895 4324
rect 2911 4380 2975 4384
rect 2911 4324 2915 4380
rect 2915 4324 2971 4380
rect 2971 4324 2975 4380
rect 2911 4320 2975 4324
rect 2991 4380 3055 4384
rect 2991 4324 2995 4380
rect 2995 4324 3051 4380
rect 3051 4324 3055 4380
rect 2991 4320 3055 4324
rect 3071 4380 3135 4384
rect 3071 4324 3075 4380
rect 3075 4324 3131 4380
rect 3131 4324 3135 4380
rect 3071 4320 3135 4324
rect 5269 4380 5333 4384
rect 5269 4324 5273 4380
rect 5273 4324 5329 4380
rect 5329 4324 5333 4380
rect 5269 4320 5333 4324
rect 5349 4380 5413 4384
rect 5349 4324 5353 4380
rect 5353 4324 5409 4380
rect 5409 4324 5413 4380
rect 5349 4320 5413 4324
rect 5429 4380 5493 4384
rect 5429 4324 5433 4380
rect 5433 4324 5489 4380
rect 5489 4324 5493 4380
rect 5429 4320 5493 4324
rect 5509 4380 5573 4384
rect 5509 4324 5513 4380
rect 5513 4324 5569 4380
rect 5569 4324 5573 4380
rect 5509 4320 5573 4324
rect 7707 4380 7771 4384
rect 7707 4324 7711 4380
rect 7711 4324 7767 4380
rect 7767 4324 7771 4380
rect 7707 4320 7771 4324
rect 7787 4380 7851 4384
rect 7787 4324 7791 4380
rect 7791 4324 7847 4380
rect 7847 4324 7851 4380
rect 7787 4320 7851 4324
rect 7867 4380 7931 4384
rect 7867 4324 7871 4380
rect 7871 4324 7927 4380
rect 7927 4324 7931 4380
rect 7867 4320 7931 4324
rect 7947 4380 8011 4384
rect 7947 4324 7951 4380
rect 7951 4324 8007 4380
rect 8007 4324 8011 4380
rect 7947 4320 8011 4324
rect 10145 4380 10209 4384
rect 10145 4324 10149 4380
rect 10149 4324 10205 4380
rect 10205 4324 10209 4380
rect 10145 4320 10209 4324
rect 10225 4380 10289 4384
rect 10225 4324 10229 4380
rect 10229 4324 10285 4380
rect 10285 4324 10289 4380
rect 10225 4320 10289 4324
rect 10305 4380 10369 4384
rect 10305 4324 10309 4380
rect 10309 4324 10365 4380
rect 10365 4324 10369 4380
rect 10305 4320 10369 4324
rect 10385 4380 10449 4384
rect 10385 4324 10389 4380
rect 10389 4324 10445 4380
rect 10445 4324 10449 4380
rect 10385 4320 10449 4324
rect 2171 3836 2235 3840
rect 2171 3780 2175 3836
rect 2175 3780 2231 3836
rect 2231 3780 2235 3836
rect 2171 3776 2235 3780
rect 2251 3836 2315 3840
rect 2251 3780 2255 3836
rect 2255 3780 2311 3836
rect 2311 3780 2315 3836
rect 2251 3776 2315 3780
rect 2331 3836 2395 3840
rect 2331 3780 2335 3836
rect 2335 3780 2391 3836
rect 2391 3780 2395 3836
rect 2331 3776 2395 3780
rect 2411 3836 2475 3840
rect 2411 3780 2415 3836
rect 2415 3780 2471 3836
rect 2471 3780 2475 3836
rect 2411 3776 2475 3780
rect 4609 3836 4673 3840
rect 4609 3780 4613 3836
rect 4613 3780 4669 3836
rect 4669 3780 4673 3836
rect 4609 3776 4673 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 7047 3836 7111 3840
rect 7047 3780 7051 3836
rect 7051 3780 7107 3836
rect 7107 3780 7111 3836
rect 7047 3776 7111 3780
rect 7127 3836 7191 3840
rect 7127 3780 7131 3836
rect 7131 3780 7187 3836
rect 7187 3780 7191 3836
rect 7127 3776 7191 3780
rect 7207 3836 7271 3840
rect 7207 3780 7211 3836
rect 7211 3780 7267 3836
rect 7267 3780 7271 3836
rect 7207 3776 7271 3780
rect 7287 3836 7351 3840
rect 7287 3780 7291 3836
rect 7291 3780 7347 3836
rect 7347 3780 7351 3836
rect 7287 3776 7351 3780
rect 9485 3836 9549 3840
rect 9485 3780 9489 3836
rect 9489 3780 9545 3836
rect 9545 3780 9549 3836
rect 9485 3776 9549 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 2831 3292 2895 3296
rect 2831 3236 2835 3292
rect 2835 3236 2891 3292
rect 2891 3236 2895 3292
rect 2831 3232 2895 3236
rect 2911 3292 2975 3296
rect 2911 3236 2915 3292
rect 2915 3236 2971 3292
rect 2971 3236 2975 3292
rect 2911 3232 2975 3236
rect 2991 3292 3055 3296
rect 2991 3236 2995 3292
rect 2995 3236 3051 3292
rect 3051 3236 3055 3292
rect 2991 3232 3055 3236
rect 3071 3292 3135 3296
rect 3071 3236 3075 3292
rect 3075 3236 3131 3292
rect 3131 3236 3135 3292
rect 3071 3232 3135 3236
rect 5269 3292 5333 3296
rect 5269 3236 5273 3292
rect 5273 3236 5329 3292
rect 5329 3236 5333 3292
rect 5269 3232 5333 3236
rect 5349 3292 5413 3296
rect 5349 3236 5353 3292
rect 5353 3236 5409 3292
rect 5409 3236 5413 3292
rect 5349 3232 5413 3236
rect 5429 3292 5493 3296
rect 5429 3236 5433 3292
rect 5433 3236 5489 3292
rect 5489 3236 5493 3292
rect 5429 3232 5493 3236
rect 5509 3292 5573 3296
rect 5509 3236 5513 3292
rect 5513 3236 5569 3292
rect 5569 3236 5573 3292
rect 5509 3232 5573 3236
rect 7707 3292 7771 3296
rect 7707 3236 7711 3292
rect 7711 3236 7767 3292
rect 7767 3236 7771 3292
rect 7707 3232 7771 3236
rect 7787 3292 7851 3296
rect 7787 3236 7791 3292
rect 7791 3236 7847 3292
rect 7847 3236 7851 3292
rect 7787 3232 7851 3236
rect 7867 3292 7931 3296
rect 7867 3236 7871 3292
rect 7871 3236 7927 3292
rect 7927 3236 7931 3292
rect 7867 3232 7931 3236
rect 7947 3292 8011 3296
rect 7947 3236 7951 3292
rect 7951 3236 8007 3292
rect 8007 3236 8011 3292
rect 7947 3232 8011 3236
rect 10145 3292 10209 3296
rect 10145 3236 10149 3292
rect 10149 3236 10205 3292
rect 10205 3236 10209 3292
rect 10145 3232 10209 3236
rect 10225 3292 10289 3296
rect 10225 3236 10229 3292
rect 10229 3236 10285 3292
rect 10285 3236 10289 3292
rect 10225 3232 10289 3236
rect 10305 3292 10369 3296
rect 10305 3236 10309 3292
rect 10309 3236 10365 3292
rect 10365 3236 10369 3292
rect 10305 3232 10369 3236
rect 10385 3292 10449 3296
rect 10385 3236 10389 3292
rect 10389 3236 10445 3292
rect 10445 3236 10449 3292
rect 10385 3232 10449 3236
rect 2171 2748 2235 2752
rect 2171 2692 2175 2748
rect 2175 2692 2231 2748
rect 2231 2692 2235 2748
rect 2171 2688 2235 2692
rect 2251 2748 2315 2752
rect 2251 2692 2255 2748
rect 2255 2692 2311 2748
rect 2311 2692 2315 2748
rect 2251 2688 2315 2692
rect 2331 2748 2395 2752
rect 2331 2692 2335 2748
rect 2335 2692 2391 2748
rect 2391 2692 2395 2748
rect 2331 2688 2395 2692
rect 2411 2748 2475 2752
rect 2411 2692 2415 2748
rect 2415 2692 2471 2748
rect 2471 2692 2475 2748
rect 2411 2688 2475 2692
rect 4609 2748 4673 2752
rect 4609 2692 4613 2748
rect 4613 2692 4669 2748
rect 4669 2692 4673 2748
rect 4609 2688 4673 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 7047 2748 7111 2752
rect 7047 2692 7051 2748
rect 7051 2692 7107 2748
rect 7107 2692 7111 2748
rect 7047 2688 7111 2692
rect 7127 2748 7191 2752
rect 7127 2692 7131 2748
rect 7131 2692 7187 2748
rect 7187 2692 7191 2748
rect 7127 2688 7191 2692
rect 7207 2748 7271 2752
rect 7207 2692 7211 2748
rect 7211 2692 7267 2748
rect 7267 2692 7271 2748
rect 7207 2688 7271 2692
rect 7287 2748 7351 2752
rect 7287 2692 7291 2748
rect 7291 2692 7347 2748
rect 7347 2692 7351 2748
rect 7287 2688 7351 2692
rect 9485 2748 9549 2752
rect 9485 2692 9489 2748
rect 9489 2692 9545 2748
rect 9545 2692 9549 2748
rect 9485 2688 9549 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 2831 2204 2895 2208
rect 2831 2148 2835 2204
rect 2835 2148 2891 2204
rect 2891 2148 2895 2204
rect 2831 2144 2895 2148
rect 2911 2204 2975 2208
rect 2911 2148 2915 2204
rect 2915 2148 2971 2204
rect 2971 2148 2975 2204
rect 2911 2144 2975 2148
rect 2991 2204 3055 2208
rect 2991 2148 2995 2204
rect 2995 2148 3051 2204
rect 3051 2148 3055 2204
rect 2991 2144 3055 2148
rect 3071 2204 3135 2208
rect 3071 2148 3075 2204
rect 3075 2148 3131 2204
rect 3131 2148 3135 2204
rect 3071 2144 3135 2148
rect 5269 2204 5333 2208
rect 5269 2148 5273 2204
rect 5273 2148 5329 2204
rect 5329 2148 5333 2204
rect 5269 2144 5333 2148
rect 5349 2204 5413 2208
rect 5349 2148 5353 2204
rect 5353 2148 5409 2204
rect 5409 2148 5413 2204
rect 5349 2144 5413 2148
rect 5429 2204 5493 2208
rect 5429 2148 5433 2204
rect 5433 2148 5489 2204
rect 5489 2148 5493 2204
rect 5429 2144 5493 2148
rect 5509 2204 5573 2208
rect 5509 2148 5513 2204
rect 5513 2148 5569 2204
rect 5569 2148 5573 2204
rect 5509 2144 5573 2148
rect 7707 2204 7771 2208
rect 7707 2148 7711 2204
rect 7711 2148 7767 2204
rect 7767 2148 7771 2204
rect 7707 2144 7771 2148
rect 7787 2204 7851 2208
rect 7787 2148 7791 2204
rect 7791 2148 7847 2204
rect 7847 2148 7851 2204
rect 7787 2144 7851 2148
rect 7867 2204 7931 2208
rect 7867 2148 7871 2204
rect 7871 2148 7927 2204
rect 7927 2148 7931 2204
rect 7867 2144 7931 2148
rect 7947 2204 8011 2208
rect 7947 2148 7951 2204
rect 7951 2148 8007 2204
rect 8007 2148 8011 2204
rect 7947 2144 8011 2148
rect 10145 2204 10209 2208
rect 10145 2148 10149 2204
rect 10149 2148 10205 2204
rect 10205 2148 10209 2204
rect 10145 2144 10209 2148
rect 10225 2204 10289 2208
rect 10225 2148 10229 2204
rect 10229 2148 10285 2204
rect 10285 2148 10289 2204
rect 10225 2144 10289 2148
rect 10305 2204 10369 2208
rect 10305 2148 10309 2204
rect 10309 2148 10365 2204
rect 10365 2148 10369 2204
rect 10305 2144 10369 2148
rect 10385 2204 10449 2208
rect 10385 2148 10389 2204
rect 10389 2148 10445 2204
rect 10445 2148 10449 2204
rect 10385 2144 10449 2148
<< metal4 >>
rect 2163 11456 2483 11472
rect 2163 11392 2171 11456
rect 2235 11392 2251 11456
rect 2315 11392 2331 11456
rect 2395 11392 2411 11456
rect 2475 11392 2483 11456
rect 2163 10382 2483 11392
rect 2163 10368 2205 10382
rect 2441 10368 2483 10382
rect 2163 10304 2171 10368
rect 2475 10304 2483 10368
rect 2163 10146 2205 10304
rect 2441 10146 2483 10304
rect 2163 9280 2483 10146
rect 2163 9216 2171 9280
rect 2235 9216 2251 9280
rect 2315 9216 2331 9280
rect 2395 9216 2411 9280
rect 2475 9216 2483 9280
rect 2163 8192 2483 9216
rect 2163 8128 2171 8192
rect 2235 8128 2251 8192
rect 2315 8128 2331 8192
rect 2395 8128 2411 8192
rect 2475 8128 2483 8192
rect 2163 8071 2483 8128
rect 2163 7835 2205 8071
rect 2441 7835 2483 8071
rect 2163 7104 2483 7835
rect 2163 7040 2171 7104
rect 2235 7040 2251 7104
rect 2315 7040 2331 7104
rect 2395 7040 2411 7104
rect 2475 7040 2483 7104
rect 2163 6016 2483 7040
rect 2163 5952 2171 6016
rect 2235 5952 2251 6016
rect 2315 5952 2331 6016
rect 2395 5952 2411 6016
rect 2475 5952 2483 6016
rect 2163 5760 2483 5952
rect 2163 5524 2205 5760
rect 2441 5524 2483 5760
rect 2163 4928 2483 5524
rect 2163 4864 2171 4928
rect 2235 4864 2251 4928
rect 2315 4864 2331 4928
rect 2395 4864 2411 4928
rect 2475 4864 2483 4928
rect 2163 3840 2483 4864
rect 2163 3776 2171 3840
rect 2235 3776 2251 3840
rect 2315 3776 2331 3840
rect 2395 3776 2411 3840
rect 2475 3776 2483 3840
rect 2163 3449 2483 3776
rect 2163 3213 2205 3449
rect 2441 3213 2483 3449
rect 2163 2752 2483 3213
rect 2163 2688 2171 2752
rect 2235 2688 2251 2752
rect 2315 2688 2331 2752
rect 2395 2688 2411 2752
rect 2475 2688 2483 2752
rect 2163 2128 2483 2688
rect 2823 11042 3143 11472
rect 2823 10912 2865 11042
rect 3101 10912 3143 11042
rect 2823 10848 2831 10912
rect 3135 10848 3143 10912
rect 2823 10806 2865 10848
rect 3101 10806 3143 10848
rect 2823 9824 3143 10806
rect 2823 9760 2831 9824
rect 2895 9760 2911 9824
rect 2975 9760 2991 9824
rect 3055 9760 3071 9824
rect 3135 9760 3143 9824
rect 2823 8736 3143 9760
rect 2823 8672 2831 8736
rect 2895 8731 2911 8736
rect 2975 8731 2991 8736
rect 3055 8731 3071 8736
rect 3135 8672 3143 8736
rect 2823 8495 2865 8672
rect 3101 8495 3143 8672
rect 2823 7648 3143 8495
rect 2823 7584 2831 7648
rect 2895 7584 2911 7648
rect 2975 7584 2991 7648
rect 3055 7584 3071 7648
rect 3135 7584 3143 7648
rect 2823 6560 3143 7584
rect 2823 6496 2831 6560
rect 2895 6496 2911 6560
rect 2975 6496 2991 6560
rect 3055 6496 3071 6560
rect 3135 6496 3143 6560
rect 2823 6420 3143 6496
rect 2823 6184 2865 6420
rect 3101 6184 3143 6420
rect 2823 5472 3143 6184
rect 2823 5408 2831 5472
rect 2895 5408 2911 5472
rect 2975 5408 2991 5472
rect 3055 5408 3071 5472
rect 3135 5408 3143 5472
rect 2823 4384 3143 5408
rect 2823 4320 2831 4384
rect 2895 4320 2911 4384
rect 2975 4320 2991 4384
rect 3055 4320 3071 4384
rect 3135 4320 3143 4384
rect 2823 4109 3143 4320
rect 2823 3873 2865 4109
rect 3101 3873 3143 4109
rect 2823 3296 3143 3873
rect 2823 3232 2831 3296
rect 2895 3232 2911 3296
rect 2975 3232 2991 3296
rect 3055 3232 3071 3296
rect 3135 3232 3143 3296
rect 2823 2208 3143 3232
rect 2823 2144 2831 2208
rect 2895 2144 2911 2208
rect 2975 2144 2991 2208
rect 3055 2144 3071 2208
rect 3135 2144 3143 2208
rect 2823 2128 3143 2144
rect 4601 11456 4921 11472
rect 4601 11392 4609 11456
rect 4673 11392 4689 11456
rect 4753 11392 4769 11456
rect 4833 11392 4849 11456
rect 4913 11392 4921 11456
rect 4601 10382 4921 11392
rect 4601 10368 4643 10382
rect 4879 10368 4921 10382
rect 4601 10304 4609 10368
rect 4913 10304 4921 10368
rect 4601 10146 4643 10304
rect 4879 10146 4921 10304
rect 4601 9280 4921 10146
rect 4601 9216 4609 9280
rect 4673 9216 4689 9280
rect 4753 9216 4769 9280
rect 4833 9216 4849 9280
rect 4913 9216 4921 9280
rect 4601 8192 4921 9216
rect 4601 8128 4609 8192
rect 4673 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4921 8192
rect 4601 8071 4921 8128
rect 4601 7835 4643 8071
rect 4879 7835 4921 8071
rect 4601 7104 4921 7835
rect 4601 7040 4609 7104
rect 4673 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4921 7104
rect 4601 6016 4921 7040
rect 4601 5952 4609 6016
rect 4673 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4921 6016
rect 4601 5760 4921 5952
rect 4601 5524 4643 5760
rect 4879 5524 4921 5760
rect 4601 4928 4921 5524
rect 4601 4864 4609 4928
rect 4673 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4921 4928
rect 4601 3840 4921 4864
rect 4601 3776 4609 3840
rect 4673 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4921 3840
rect 4601 3449 4921 3776
rect 4601 3213 4643 3449
rect 4879 3213 4921 3449
rect 4601 2752 4921 3213
rect 4601 2688 4609 2752
rect 4673 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4921 2752
rect 4601 2128 4921 2688
rect 5261 11042 5581 11472
rect 5261 10912 5303 11042
rect 5539 10912 5581 11042
rect 5261 10848 5269 10912
rect 5573 10848 5581 10912
rect 5261 10806 5303 10848
rect 5539 10806 5581 10848
rect 5261 9824 5581 10806
rect 5261 9760 5269 9824
rect 5333 9760 5349 9824
rect 5413 9760 5429 9824
rect 5493 9760 5509 9824
rect 5573 9760 5581 9824
rect 5261 8736 5581 9760
rect 5261 8672 5269 8736
rect 5333 8731 5349 8736
rect 5413 8731 5429 8736
rect 5493 8731 5509 8736
rect 5573 8672 5581 8736
rect 5261 8495 5303 8672
rect 5539 8495 5581 8672
rect 5261 7648 5581 8495
rect 5261 7584 5269 7648
rect 5333 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5581 7648
rect 5261 6560 5581 7584
rect 5261 6496 5269 6560
rect 5333 6496 5349 6560
rect 5413 6496 5429 6560
rect 5493 6496 5509 6560
rect 5573 6496 5581 6560
rect 5261 6420 5581 6496
rect 5261 6184 5303 6420
rect 5539 6184 5581 6420
rect 5261 5472 5581 6184
rect 5261 5408 5269 5472
rect 5333 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5581 5472
rect 5261 4384 5581 5408
rect 5261 4320 5269 4384
rect 5333 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5581 4384
rect 5261 4109 5581 4320
rect 5261 3873 5303 4109
rect 5539 3873 5581 4109
rect 5261 3296 5581 3873
rect 5261 3232 5269 3296
rect 5333 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5581 3296
rect 5261 2208 5581 3232
rect 5261 2144 5269 2208
rect 5333 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5581 2208
rect 5261 2128 5581 2144
rect 7039 11456 7359 11472
rect 7039 11392 7047 11456
rect 7111 11392 7127 11456
rect 7191 11392 7207 11456
rect 7271 11392 7287 11456
rect 7351 11392 7359 11456
rect 7039 10382 7359 11392
rect 7039 10368 7081 10382
rect 7317 10368 7359 10382
rect 7039 10304 7047 10368
rect 7351 10304 7359 10368
rect 7039 10146 7081 10304
rect 7317 10146 7359 10304
rect 7039 9280 7359 10146
rect 7039 9216 7047 9280
rect 7111 9216 7127 9280
rect 7191 9216 7207 9280
rect 7271 9216 7287 9280
rect 7351 9216 7359 9280
rect 7039 8192 7359 9216
rect 7039 8128 7047 8192
rect 7111 8128 7127 8192
rect 7191 8128 7207 8192
rect 7271 8128 7287 8192
rect 7351 8128 7359 8192
rect 7039 8071 7359 8128
rect 7039 7835 7081 8071
rect 7317 7835 7359 8071
rect 7039 7104 7359 7835
rect 7039 7040 7047 7104
rect 7111 7040 7127 7104
rect 7191 7040 7207 7104
rect 7271 7040 7287 7104
rect 7351 7040 7359 7104
rect 7039 6016 7359 7040
rect 7039 5952 7047 6016
rect 7111 5952 7127 6016
rect 7191 5952 7207 6016
rect 7271 5952 7287 6016
rect 7351 5952 7359 6016
rect 7039 5760 7359 5952
rect 7039 5524 7081 5760
rect 7317 5524 7359 5760
rect 7039 4928 7359 5524
rect 7039 4864 7047 4928
rect 7111 4864 7127 4928
rect 7191 4864 7207 4928
rect 7271 4864 7287 4928
rect 7351 4864 7359 4928
rect 7039 3840 7359 4864
rect 7039 3776 7047 3840
rect 7111 3776 7127 3840
rect 7191 3776 7207 3840
rect 7271 3776 7287 3840
rect 7351 3776 7359 3840
rect 7039 3449 7359 3776
rect 7039 3213 7081 3449
rect 7317 3213 7359 3449
rect 7039 2752 7359 3213
rect 7039 2688 7047 2752
rect 7111 2688 7127 2752
rect 7191 2688 7207 2752
rect 7271 2688 7287 2752
rect 7351 2688 7359 2752
rect 7039 2128 7359 2688
rect 7699 11042 8019 11472
rect 7699 10912 7741 11042
rect 7977 10912 8019 11042
rect 7699 10848 7707 10912
rect 8011 10848 8019 10912
rect 7699 10806 7741 10848
rect 7977 10806 8019 10848
rect 7699 9824 8019 10806
rect 7699 9760 7707 9824
rect 7771 9760 7787 9824
rect 7851 9760 7867 9824
rect 7931 9760 7947 9824
rect 8011 9760 8019 9824
rect 7699 8736 8019 9760
rect 7699 8672 7707 8736
rect 7771 8731 7787 8736
rect 7851 8731 7867 8736
rect 7931 8731 7947 8736
rect 8011 8672 8019 8736
rect 7699 8495 7741 8672
rect 7977 8495 8019 8672
rect 7699 7648 8019 8495
rect 7699 7584 7707 7648
rect 7771 7584 7787 7648
rect 7851 7584 7867 7648
rect 7931 7584 7947 7648
rect 8011 7584 8019 7648
rect 7699 6560 8019 7584
rect 7699 6496 7707 6560
rect 7771 6496 7787 6560
rect 7851 6496 7867 6560
rect 7931 6496 7947 6560
rect 8011 6496 8019 6560
rect 7699 6420 8019 6496
rect 7699 6184 7741 6420
rect 7977 6184 8019 6420
rect 7699 5472 8019 6184
rect 7699 5408 7707 5472
rect 7771 5408 7787 5472
rect 7851 5408 7867 5472
rect 7931 5408 7947 5472
rect 8011 5408 8019 5472
rect 7699 4384 8019 5408
rect 7699 4320 7707 4384
rect 7771 4320 7787 4384
rect 7851 4320 7867 4384
rect 7931 4320 7947 4384
rect 8011 4320 8019 4384
rect 7699 4109 8019 4320
rect 7699 3873 7741 4109
rect 7977 3873 8019 4109
rect 7699 3296 8019 3873
rect 7699 3232 7707 3296
rect 7771 3232 7787 3296
rect 7851 3232 7867 3296
rect 7931 3232 7947 3296
rect 8011 3232 8019 3296
rect 7699 2208 8019 3232
rect 7699 2144 7707 2208
rect 7771 2144 7787 2208
rect 7851 2144 7867 2208
rect 7931 2144 7947 2208
rect 8011 2144 8019 2208
rect 7699 2128 8019 2144
rect 9477 11456 9797 11472
rect 9477 11392 9485 11456
rect 9549 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9797 11456
rect 9477 10382 9797 11392
rect 9477 10368 9519 10382
rect 9755 10368 9797 10382
rect 9477 10304 9485 10368
rect 9789 10304 9797 10368
rect 9477 10146 9519 10304
rect 9755 10146 9797 10304
rect 9477 9280 9797 10146
rect 9477 9216 9485 9280
rect 9549 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9797 9280
rect 9477 8192 9797 9216
rect 9477 8128 9485 8192
rect 9549 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9797 8192
rect 9477 8071 9797 8128
rect 9477 7835 9519 8071
rect 9755 7835 9797 8071
rect 9477 7104 9797 7835
rect 9477 7040 9485 7104
rect 9549 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9797 7104
rect 9477 6016 9797 7040
rect 9477 5952 9485 6016
rect 9549 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9797 6016
rect 9477 5760 9797 5952
rect 9477 5524 9519 5760
rect 9755 5524 9797 5760
rect 9477 4928 9797 5524
rect 9477 4864 9485 4928
rect 9549 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9797 4928
rect 9477 3840 9797 4864
rect 9477 3776 9485 3840
rect 9549 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9797 3840
rect 9477 3449 9797 3776
rect 9477 3213 9519 3449
rect 9755 3213 9797 3449
rect 9477 2752 9797 3213
rect 9477 2688 9485 2752
rect 9549 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9797 2752
rect 9477 2128 9797 2688
rect 10137 11042 10457 11472
rect 10137 10912 10179 11042
rect 10415 10912 10457 11042
rect 10137 10848 10145 10912
rect 10449 10848 10457 10912
rect 10137 10806 10179 10848
rect 10415 10806 10457 10848
rect 10137 9824 10457 10806
rect 10137 9760 10145 9824
rect 10209 9760 10225 9824
rect 10289 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10457 9824
rect 10137 8736 10457 9760
rect 10137 8672 10145 8736
rect 10209 8731 10225 8736
rect 10289 8731 10305 8736
rect 10369 8731 10385 8736
rect 10449 8672 10457 8736
rect 10137 8495 10179 8672
rect 10415 8495 10457 8672
rect 10137 7648 10457 8495
rect 10137 7584 10145 7648
rect 10209 7584 10225 7648
rect 10289 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10457 7648
rect 10137 6560 10457 7584
rect 10137 6496 10145 6560
rect 10209 6496 10225 6560
rect 10289 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10457 6560
rect 10137 6420 10457 6496
rect 10137 6184 10179 6420
rect 10415 6184 10457 6420
rect 10137 5472 10457 6184
rect 10137 5408 10145 5472
rect 10209 5408 10225 5472
rect 10289 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10457 5472
rect 10137 4384 10457 5408
rect 10137 4320 10145 4384
rect 10209 4320 10225 4384
rect 10289 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10457 4384
rect 10137 4109 10457 4320
rect 10137 3873 10179 4109
rect 10415 3873 10457 4109
rect 10137 3296 10457 3873
rect 10137 3232 10145 3296
rect 10209 3232 10225 3296
rect 10289 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10457 3296
rect 10137 2208 10457 3232
rect 10137 2144 10145 2208
rect 10209 2144 10225 2208
rect 10289 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10457 2208
rect 10137 2128 10457 2144
<< via4 >>
rect 2205 10368 2441 10382
rect 2205 10304 2235 10368
rect 2235 10304 2251 10368
rect 2251 10304 2315 10368
rect 2315 10304 2331 10368
rect 2331 10304 2395 10368
rect 2395 10304 2411 10368
rect 2411 10304 2441 10368
rect 2205 10146 2441 10304
rect 2205 7835 2441 8071
rect 2205 5524 2441 5760
rect 2205 3213 2441 3449
rect 2865 10912 3101 11042
rect 2865 10848 2895 10912
rect 2895 10848 2911 10912
rect 2911 10848 2975 10912
rect 2975 10848 2991 10912
rect 2991 10848 3055 10912
rect 3055 10848 3071 10912
rect 3071 10848 3101 10912
rect 2865 10806 3101 10848
rect 2865 8672 2895 8731
rect 2895 8672 2911 8731
rect 2911 8672 2975 8731
rect 2975 8672 2991 8731
rect 2991 8672 3055 8731
rect 3055 8672 3071 8731
rect 3071 8672 3101 8731
rect 2865 8495 3101 8672
rect 2865 6184 3101 6420
rect 2865 3873 3101 4109
rect 4643 10368 4879 10382
rect 4643 10304 4673 10368
rect 4673 10304 4689 10368
rect 4689 10304 4753 10368
rect 4753 10304 4769 10368
rect 4769 10304 4833 10368
rect 4833 10304 4849 10368
rect 4849 10304 4879 10368
rect 4643 10146 4879 10304
rect 4643 7835 4879 8071
rect 4643 5524 4879 5760
rect 4643 3213 4879 3449
rect 5303 10912 5539 11042
rect 5303 10848 5333 10912
rect 5333 10848 5349 10912
rect 5349 10848 5413 10912
rect 5413 10848 5429 10912
rect 5429 10848 5493 10912
rect 5493 10848 5509 10912
rect 5509 10848 5539 10912
rect 5303 10806 5539 10848
rect 5303 8672 5333 8731
rect 5333 8672 5349 8731
rect 5349 8672 5413 8731
rect 5413 8672 5429 8731
rect 5429 8672 5493 8731
rect 5493 8672 5509 8731
rect 5509 8672 5539 8731
rect 5303 8495 5539 8672
rect 5303 6184 5539 6420
rect 5303 3873 5539 4109
rect 7081 10368 7317 10382
rect 7081 10304 7111 10368
rect 7111 10304 7127 10368
rect 7127 10304 7191 10368
rect 7191 10304 7207 10368
rect 7207 10304 7271 10368
rect 7271 10304 7287 10368
rect 7287 10304 7317 10368
rect 7081 10146 7317 10304
rect 7081 7835 7317 8071
rect 7081 5524 7317 5760
rect 7081 3213 7317 3449
rect 7741 10912 7977 11042
rect 7741 10848 7771 10912
rect 7771 10848 7787 10912
rect 7787 10848 7851 10912
rect 7851 10848 7867 10912
rect 7867 10848 7931 10912
rect 7931 10848 7947 10912
rect 7947 10848 7977 10912
rect 7741 10806 7977 10848
rect 7741 8672 7771 8731
rect 7771 8672 7787 8731
rect 7787 8672 7851 8731
rect 7851 8672 7867 8731
rect 7867 8672 7931 8731
rect 7931 8672 7947 8731
rect 7947 8672 7977 8731
rect 7741 8495 7977 8672
rect 7741 6184 7977 6420
rect 7741 3873 7977 4109
rect 9519 10368 9755 10382
rect 9519 10304 9549 10368
rect 9549 10304 9565 10368
rect 9565 10304 9629 10368
rect 9629 10304 9645 10368
rect 9645 10304 9709 10368
rect 9709 10304 9725 10368
rect 9725 10304 9755 10368
rect 9519 10146 9755 10304
rect 9519 7835 9755 8071
rect 9519 5524 9755 5760
rect 9519 3213 9755 3449
rect 10179 10912 10415 11042
rect 10179 10848 10209 10912
rect 10209 10848 10225 10912
rect 10225 10848 10289 10912
rect 10289 10848 10305 10912
rect 10305 10848 10369 10912
rect 10369 10848 10385 10912
rect 10385 10848 10415 10912
rect 10179 10806 10415 10848
rect 10179 8672 10209 8731
rect 10209 8672 10225 8731
rect 10225 8672 10289 8731
rect 10289 8672 10305 8731
rect 10305 8672 10369 8731
rect 10369 8672 10385 8731
rect 10385 8672 10415 8731
rect 10179 8495 10415 8672
rect 10179 6184 10415 6420
rect 10179 3873 10415 4109
<< metal5 >>
rect 1056 11042 10904 11084
rect 1056 10806 2865 11042
rect 3101 10806 5303 11042
rect 5539 10806 7741 11042
rect 7977 10806 10179 11042
rect 10415 10806 10904 11042
rect 1056 10764 10904 10806
rect 1056 10382 10904 10424
rect 1056 10146 2205 10382
rect 2441 10146 4643 10382
rect 4879 10146 7081 10382
rect 7317 10146 9519 10382
rect 9755 10146 10904 10382
rect 1056 10104 10904 10146
rect 1056 8731 10904 8773
rect 1056 8495 2865 8731
rect 3101 8495 5303 8731
rect 5539 8495 7741 8731
rect 7977 8495 10179 8731
rect 10415 8495 10904 8731
rect 1056 8453 10904 8495
rect 1056 8071 10904 8113
rect 1056 7835 2205 8071
rect 2441 7835 4643 8071
rect 4879 7835 7081 8071
rect 7317 7835 9519 8071
rect 9755 7835 10904 8071
rect 1056 7793 10904 7835
rect 1056 6420 10904 6462
rect 1056 6184 2865 6420
rect 3101 6184 5303 6420
rect 5539 6184 7741 6420
rect 7977 6184 10179 6420
rect 10415 6184 10904 6420
rect 1056 6142 10904 6184
rect 1056 5760 10904 5802
rect 1056 5524 2205 5760
rect 2441 5524 4643 5760
rect 4879 5524 7081 5760
rect 7317 5524 9519 5760
rect 9755 5524 10904 5760
rect 1056 5482 10904 5524
rect 1056 4109 10904 4151
rect 1056 3873 2865 4109
rect 3101 3873 5303 4109
rect 5539 3873 7741 4109
rect 7977 3873 10179 4109
rect 10415 3873 10904 4109
rect 1056 3831 10904 3873
rect 1056 3449 10904 3491
rect 1056 3213 2205 3449
rect 2441 3213 4643 3449
rect 4879 3213 7081 3449
rect 7317 3213 9519 3449
rect 9755 3213 10904 3449
rect 1056 3171 10904 3213
use sky130_fd_sc_hd__nor2_4  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6072 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10028 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9016 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _114_
timestamp 1704896540
transform 1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_4  _115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_4  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 1704896540
transform -1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 1704896540
transform -1 0 8372 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _120_
timestamp 1704896540
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _121_
timestamp 1704896540
transform -1 0 7912 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1704896540
transform 1 0 8372 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _123_
timestamp 1704896540
transform 1 0 5796 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _128_
timestamp 1704896540
transform 1 0 9108 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10212 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _130_
timestamp 1704896540
transform 1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _131_
timestamp 1704896540
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _132_
timestamp 1704896540
transform -1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _133_
timestamp 1704896540
transform -1 0 10212 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _134_
timestamp 1704896540
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _137_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1704896540
transform -1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _140_
timestamp 1704896540
transform 1 0 7820 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 1704896540
transform -1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _143_
timestamp 1704896540
transform -1 0 9752 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1704896540
transform 1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _145_
timestamp 1704896540
transform -1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10212 0 1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_2  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8464 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _148_
timestamp 1704896540
transform -1 0 6256 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _149_
timestamp 1704896540
transform -1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _150_
timestamp 1704896540
transform -1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _151_
timestamp 1704896540
transform 1 0 6900 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _152_
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1704896540
transform -1 0 7176 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _154_
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _155_
timestamp 1704896540
transform -1 0 8648 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _156_
timestamp 1704896540
transform 1 0 7360 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _157_
timestamp 1704896540
transform -1 0 7820 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _158_
timestamp 1704896540
transform -1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5336 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _160_
timestamp 1704896540
transform 1 0 3956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _163_
timestamp 1704896540
transform -1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _164_
timestamp 1704896540
transform -1 0 3680 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _165_
timestamp 1704896540
transform 1 0 2208 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _166_
timestamp 1704896540
transform -1 0 2484 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _167_
timestamp 1704896540
transform 1 0 1472 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1704896540
transform 1 0 3864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4324 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1704896540
transform -1 0 5244 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4324 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1704896540
transform 1 0 4508 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 1704896540
transform -1 0 4508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4784 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _176_
timestamp 1704896540
transform -1 0 2668 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _177_
timestamp 1704896540
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _178_
timestamp 1704896540
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _179_
timestamp 1704896540
transform -1 0 3220 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _180_
timestamp 1704896540
transform 1 0 2116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _181_
timestamp 1704896540
transform -1 0 2484 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _182_
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _184_
timestamp 1704896540
transform 1 0 4968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _185_
timestamp 1704896540
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _186_
timestamp 1704896540
transform 1 0 4140 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _187_
timestamp 1704896540
transform 1 0 4232 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _188_
timestamp 1704896540
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _189_
timestamp 1704896540
transform -1 0 2760 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _190_
timestamp 1704896540
transform -1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 1704896540
transform -1 0 3772 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _192_
timestamp 1704896540
transform 1 0 3220 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _193_
timestamp 1704896540
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _194_
timestamp 1704896540
transform -1 0 2484 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _195_
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1704896540
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _197_
timestamp 1704896540
transform -1 0 4324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _198_
timestamp 1704896540
transform -1 0 5796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _199_
timestamp 1704896540
transform 1 0 4140 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _200_
timestamp 1704896540
transform 1 0 4324 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _201_
timestamp 1704896540
transform -1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _202_
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _204_
timestamp 1704896540
transform -1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _205_
timestamp 1704896540
transform -1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _206_
timestamp 1704896540
transform -1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _207_
timestamp 1704896540
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _209_
timestamp 1704896540
transform 1 0 2300 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _210_
timestamp 1704896540
transform 1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1704896540
transform -1 0 4968 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _214_
timestamp 1704896540
transform -1 0 8832 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _215_
timestamp 1704896540
transform 1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _216_
timestamp 1704896540
transform -1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7544 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7544 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1704896540
transform -1 0 6716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1704896540
transform -1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1704896540
transform -1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1704896540
transform 1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1704896540
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1704896540
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1704896540
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_70
timestamp 1704896540
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_90
timestamp 1704896540
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1704896540
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_13
timestamp 1704896540
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_17
timestamp 1704896540
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_24
timestamp 1704896540
transform 1 0 3312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_30
timestamp 1704896540
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_35
timestamp 1704896540
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1704896540
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_76
timestamp 1704896540
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_86
timestamp 1704896540
transform 1 0 9016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 1704896540
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_12
timestamp 1704896540
transform 1 0 2208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_54
timestamp 1704896540
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_60
timestamp 1704896540
transform 1 0 6624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_76
timestamp 1704896540
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_33
timestamp 1704896540
transform 1 0 4140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_37
timestamp 1704896540
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_63
timestamp 1704896540
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_78
timestamp 1704896540
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_97
timestamp 1704896540
transform 1 0 10028 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1704896540
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1704896540
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_49
timestamp 1704896540
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_65
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_92
timestamp 1704896540
transform 1 0 9568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_100
timestamp 1704896540
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_10
timestamp 1704896540
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_18
timestamp 1704896540
transform 1 0 2760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_33
timestamp 1704896540
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_74
timestamp 1704896540
transform 1 0 7912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_97
timestamp 1704896540
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_51
timestamp 1704896540
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_67
timestamp 1704896540
transform 1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_99
timestamp 1704896540
transform 1 0 10212 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_6
timestamp 1704896540
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_38
timestamp 1704896540
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_49
timestamp 1704896540
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_68
timestamp 1704896540
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1704896540
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_102
timestamp 1704896540
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_6
timestamp 1704896540
transform 1 0 1656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_10
timestamp 1704896540
transform 1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_17
timestamp 1704896540
transform 1 0 2668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_23
timestamp 1704896540
transform 1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_42
timestamp 1704896540
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_50
timestamp 1704896540
transform 1 0 5704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_73
timestamp 1704896540
transform 1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_88
timestamp 1704896540
transform 1 0 9200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_22
timestamp 1704896540
transform 1 0 3128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_32
timestamp 1704896540
transform 1 0 4048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_49
timestamp 1704896540
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_64
timestamp 1704896540
transform 1 0 6992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_80
timestamp 1704896540
transform 1 0 8464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_7
timestamp 1704896540
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1704896540
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_30
timestamp 1704896540
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_40
timestamp 1704896540
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1704896540
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1704896540
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1704896540
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1704896540
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_99
timestamp 1704896540
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_9
timestamp 1704896540
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_15
timestamp 1704896540
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_21
timestamp 1704896540
transform 1 0 3036 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_31
timestamp 1704896540
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_44
timestamp 1704896540
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_65
timestamp 1704896540
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_79
timestamp 1704896540
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_91
timestamp 1704896540
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_20
timestamp 1704896540
transform 1 0 2944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_49
timestamp 1704896540
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_61
timestamp 1704896540
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1704896540
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_7
timestamp 1704896540
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_11
timestamp 1704896540
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_19
timestamp 1704896540
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_46
timestamp 1704896540
transform 1 0 5336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_66
timestamp 1704896540
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_83
timestamp 1704896540
transform 1 0 8740 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_95
timestamp 1704896540
transform 1 0 9844 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_34
timestamp 1704896540
transform 1 0 4232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_50
timestamp 1704896540
transform 1 0 5704 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_63
timestamp 1704896540
transform 1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1704896540
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_88
timestamp 1704896540
transform 1 0 9200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_100
timestamp 1704896540
transform 1 0 10304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 10580 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform -1 0 8740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform -1 0 5704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1704896540
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1704896540
transform -1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1704896540
transform -1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1704896540
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1704896540
transform -1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1704896540
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1704896540
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1704896540
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10580 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input20
timestamp 1704896540
transform -1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output21
timestamp 1704896540
transform -1 0 5612 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1704896540
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1704896540
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1704896540
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output29
timestamp 1704896540
transform -1 0 2208 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_17
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_18
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_19
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_20
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_22
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_26
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_27
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_28
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_29
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_30
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_31
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_32
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_33
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer1
timestamp 1704896540
transform -1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5428 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 1704896540
transform 1 0 8004 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7084 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer5
timestamp 1704896540
transform 1 0 8648 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer6
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 1704896540
transform -1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer8
timestamp 1704896540
transform -1 0 5336 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 1704896540
transform -1 0 5336 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer10
timestamp 1704896540
transform 1 0 9660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer11
timestamp 1704896540
transform -1 0 10212 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer12
timestamp 1704896540
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer13
timestamp 1704896540
transform 1 0 7268 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_41
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_42
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_43
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_44
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_45
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_46
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_47
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_48
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_49
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_50
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_51
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_52
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_53
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_54
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_55
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_56
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_57
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_59
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_60
timestamp 1704896540
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 2823 2128 3143 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5261 2128 5581 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7699 2128 8019 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10137 2128 10457 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3831 10904 4151 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6142 10904 6462 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8453 10904 8773 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10764 10904 11084 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2163 2128 2483 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4601 2128 4921 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7039 2128 7359 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9477 2128 9797 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3171 10904 3491 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5482 10904 5802 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7793 10904 8113 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 10104 10904 10424 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 a[0]
port 2 nsew signal input
flabel metal3 s 11198 4768 11998 4888 0 FreeSans 480 0 0 0 a[1]
port 3 nsew signal input
flabel metal3 s 11198 8848 11998 8968 0 FreeSans 480 0 0 0 a[2]
port 4 nsew signal input
flabel metal2 s 7746 13342 7802 14142 0 FreeSans 224 90 0 0 a[3]
port 5 nsew signal input
flabel metal2 s 4526 13342 4582 14142 0 FreeSans 224 90 0 0 a[4]
port 6 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 a[5]
port 7 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 a[6]
port 8 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 a[7]
port 9 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 b[0]
port 10 nsew signal input
flabel metal3 s 11198 5448 11998 5568 0 FreeSans 480 0 0 0 b[1]
port 11 nsew signal input
flabel metal3 s 11198 8168 11998 8288 0 FreeSans 480 0 0 0 b[2]
port 12 nsew signal input
flabel metal2 s 7102 13342 7158 14142 0 FreeSans 224 90 0 0 b[3]
port 13 nsew signal input
flabel metal2 s 3882 13342 3938 14142 0 FreeSans 224 90 0 0 b[4]
port 14 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 b[5]
port 15 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 b[6]
port 16 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 b[7]
port 17 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 cin
port 18 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 cout
port 19 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 op[0]
port 20 nsew signal input
flabel metal3 s 11198 6808 11998 6928 0 FreeSans 480 0 0 0 op[1]
port 21 nsew signal input
flabel metal3 s 11198 6128 11998 6248 0 FreeSans 480 0 0 0 op[2]
port 22 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 result[0]
port 23 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 result[1]
port 24 nsew signal output
flabel metal3 s 11198 7488 11998 7608 0 FreeSans 480 0 0 0 result[2]
port 25 nsew signal output
flabel metal2 s 5814 13342 5870 14142 0 FreeSans 224 90 0 0 result[3]
port 26 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 result[4]
port 27 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 result[5]
port 28 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 result[6]
port 29 nsew signal output
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 result[7]
port 30 nsew signal output
rlabel metal1 5980 10880 5980 10880 0 VGND
rlabel metal1 5980 11424 5980 11424 0 VPWR
rlabel metal2 2622 7956 2622 7956 0 _000_
rlabel metal1 2162 7514 2162 7514 0 _001_
rlabel metal2 1610 8092 1610 8092 0 _002_
rlabel metal1 2484 7854 2484 7854 0 _003_
rlabel metal1 3496 7922 3496 7922 0 _004_
rlabel metal1 2047 7786 2047 7786 0 _005_
rlabel metal2 2070 8092 2070 8092 0 _006_
rlabel metal1 5290 7820 5290 7820 0 _007_
rlabel metal1 4416 6086 4416 6086 0 _008_
rlabel metal1 4738 7956 4738 7956 0 _009_
rlabel metal2 4186 7038 4186 7038 0 _010_
rlabel metal1 4922 5338 4922 5338 0 _011_
rlabel metal1 3174 5746 3174 5746 0 _012_
rlabel metal1 2024 5338 2024 5338 0 _013_
rlabel metal1 1932 5678 1932 5678 0 _014_
rlabel metal1 2438 6392 2438 6392 0 _015_
rlabel metal1 3404 5542 3404 5542 0 _016_
rlabel metal1 2047 5610 2047 5610 0 _017_
rlabel metal2 2070 5916 2070 5916 0 _018_
rlabel metal2 5474 5882 5474 5882 0 _019_
rlabel metal1 5566 5644 5566 5644 0 _020_
rlabel metal1 5612 3910 5612 3910 0 _021_
rlabel metal1 4738 5678 4738 5678 0 _022_
rlabel metal2 5750 4998 5750 4998 0 _023_
rlabel metal1 4646 3026 4646 3026 0 _024_
rlabel metal1 5106 3060 5106 3060 0 _025_
rlabel metal1 5060 3570 5060 3570 0 _026_
rlabel metal1 3726 3162 3726 3162 0 _027_
rlabel metal1 4538 3094 4538 3094 0 _028_
rlabel metal1 3818 3434 3818 3434 0 _029_
rlabel metal1 3128 3026 3128 3026 0 _030_
rlabel metal2 2714 3264 2714 3264 0 _031_
rlabel metal1 5750 3570 5750 3570 0 _032_
rlabel metal2 4554 3332 4554 3332 0 _033_
rlabel metal1 5060 3366 5060 3366 0 _034_
rlabel metal1 7866 3536 7866 3536 0 _035_
rlabel metal2 7038 3264 7038 3264 0 _036_
rlabel metal1 7636 3162 7636 3162 0 _037_
rlabel metal1 7544 3638 7544 3638 0 _038_
rlabel metal2 1794 4590 1794 4590 0 _039_
rlabel metal1 8648 3026 8648 3026 0 _040_
rlabel metal1 9568 3026 9568 3026 0 _041_
rlabel metal1 8878 3162 8878 3162 0 _042_
rlabel metal1 5612 7854 5612 7854 0 _043_
rlabel metal1 9246 3162 9246 3162 0 _044_
rlabel metal1 9798 3162 9798 3162 0 _045_
rlabel metal1 2346 5644 2346 5644 0 _046_
rlabel metal1 8372 6698 8372 6698 0 _047_
rlabel metal1 8786 4046 8786 4046 0 _048_
rlabel metal1 8372 5202 8372 5202 0 _049_
rlabel metal1 9108 5066 9108 5066 0 _050_
rlabel metal1 7820 4794 7820 4794 0 _051_
rlabel metal1 6762 5712 6762 5712 0 _052_
rlabel metal2 2254 6596 2254 6596 0 _053_
rlabel metal1 8050 5270 8050 5270 0 _054_
rlabel metal2 7498 5474 7498 5474 0 _055_
rlabel metal2 8786 5304 8786 5304 0 _056_
rlabel metal1 6762 7480 6762 7480 0 _057_
rlabel metal1 6946 7242 6946 7242 0 _058_
rlabel metal1 3082 9962 3082 9962 0 _059_
rlabel metal1 6992 5338 6992 5338 0 _060_
rlabel metal1 9522 5678 9522 5678 0 _061_
rlabel metal1 10074 6766 10074 6766 0 _062_
rlabel metal1 8878 4590 8878 4590 0 _063_
rlabel metal2 9154 6596 9154 6596 0 _064_
rlabel metal1 9338 7242 9338 7242 0 _065_
rlabel metal2 8602 8092 8602 8092 0 _066_
rlabel metal2 8878 7582 8878 7582 0 _067_
rlabel metal1 8786 7344 8786 7344 0 _068_
rlabel metal1 8786 6970 8786 6970 0 _069_
rlabel metal1 7958 7310 7958 7310 0 _070_
rlabel metal1 7544 7514 7544 7514 0 _071_
rlabel metal1 8326 7956 8326 7956 0 _072_
rlabel metal2 7130 7548 7130 7548 0 _073_
rlabel metal1 9108 8398 9108 8398 0 _074_
rlabel metal1 9430 8602 9430 8602 0 _075_
rlabel metal1 10212 6834 10212 6834 0 _076_
rlabel metal1 9522 8058 9522 8058 0 _077_
rlabel metal2 8602 9588 8602 9588 0 _078_
rlabel metal1 7406 10778 7406 10778 0 _079_
rlabel metal1 6302 10064 6302 10064 0 _080_
rlabel metal2 6210 10234 6210 10234 0 _081_
rlabel metal1 7590 9486 7590 9486 0 _082_
rlabel metal2 7038 9758 7038 9758 0 _083_
rlabel metal1 6440 9690 6440 9690 0 _084_
rlabel metal2 6670 10268 6670 10268 0 _085_
rlabel metal1 8050 9962 8050 9962 0 _086_
rlabel metal1 5244 9962 5244 9962 0 _087_
rlabel metal1 7866 9588 7866 9588 0 _088_
rlabel metal1 5474 9928 5474 9928 0 _089_
rlabel metal2 2714 9792 2714 9792 0 _090_
rlabel metal1 3128 9554 3128 9554 0 _091_
rlabel metal1 2208 9418 2208 9418 0 _092_
rlabel metal2 1702 10234 1702 10234 0 _093_
rlabel metal2 2530 9826 2530 9826 0 _094_
rlabel metal1 3726 10098 3726 10098 0 _095_
rlabel metal1 2139 9962 2139 9962 0 _096_
rlabel metal1 2116 9690 2116 9690 0 _097_
rlabel metal1 4186 10030 4186 10030 0 _098_
rlabel metal2 4462 10234 4462 10234 0 _099_
rlabel metal1 4186 7514 4186 7514 0 _100_
rlabel metal1 4876 9554 4876 9554 0 _101_
rlabel metal1 4892 7446 4892 7446 0 _102_
rlabel metal1 4738 7242 4738 7242 0 _103_
rlabel metal2 5198 7684 5198 7684 0 _104_
rlabel metal2 8418 1588 8418 1588 0 a[0]
rlabel metal2 10534 5015 10534 5015 0 a[1]
rlabel via2 10534 8925 10534 8925 0 a[2]
rlabel metal2 8004 13396 8004 13396 0 a[3]
rlabel metal1 5106 11186 5106 11186 0 a[4]
rlabel metal3 751 8908 751 8908 0 a[5]
rlabel metal3 751 6188 751 6188 0 a[6]
rlabel metal2 4554 1588 4554 1588 0 a[7]
rlabel metal2 7590 3196 7590 3196 0 alu0.result
rlabel metal2 6486 5372 6486 5372 0 alu1.result
rlabel metal2 6578 7684 6578 7684 0 alu2.result
rlabel metal1 5796 10234 5796 10234 0 alu3.result
rlabel metal1 1794 10234 1794 10234 0 alu4.result
rlabel metal1 1794 7378 1794 7378 0 alu5.result
rlabel metal1 1978 5236 1978 5236 0 alu6.result
rlabel metal2 2254 3196 2254 3196 0 alu7.result
rlabel metal2 9706 1588 9706 1588 0 b[0]
rlabel metal1 10580 5678 10580 5678 0 b[1]
rlabel metal2 10534 8041 10534 8041 0 b[2]
rlabel metal1 7682 11866 7682 11866 0 b[3]
rlabel metal1 4048 11118 4048 11118 0 b[4]
rlabel metal3 751 7548 751 7548 0 b[5]
rlabel metal3 751 4828 751 4828 0 b[6]
rlabel metal2 3910 1588 3910 1588 0 b[7]
rlabel metal2 9062 1588 9062 1588 0 cin
rlabel metal2 5198 1554 5198 1554 0 cout
rlabel metal1 8970 2618 8970 2618 0 net1
rlabel metal1 10166 5780 10166 5780 0 net10
rlabel metal1 10028 8466 10028 8466 0 net11
rlabel metal2 8326 10268 8326 10268 0 net12
rlabel metal2 3910 10506 3910 10506 0 net13
rlabel metal1 2024 7446 2024 7446 0 net14
rlabel metal1 3174 5610 3174 5610 0 net15
rlabel metal1 4094 2958 4094 2958 0 net16
rlabel metal2 9338 2689 9338 2689 0 net17
rlabel metal1 6624 2618 6624 2618 0 net18
rlabel metal1 7866 6766 7866 6766 0 net19
rlabel metal1 9706 5202 9706 5202 0 net2
rlabel metal2 6762 6562 6762 6562 0 net20
rlabel metal1 5612 2414 5612 2414 0 net21
rlabel metal1 7820 2822 7820 2822 0 net22
rlabel metal1 7084 2414 7084 2414 0 net23
rlabel metal1 8050 8058 8050 8058 0 net24
rlabel metal1 6118 10778 6118 10778 0 net25
rlabel metal1 1794 10642 1794 10642 0 net26
rlabel metal1 1748 7514 1748 7514 0 net27
rlabel metal1 1748 5202 1748 5202 0 net28
rlabel metal2 2070 3332 2070 3332 0 net29
rlabel metal2 9982 8670 9982 8670 0 net3
rlabel metal2 5290 10438 5290 10438 0 net30
rlabel metal2 4278 10812 4278 10812 0 net31
rlabel metal1 7130 11220 7130 11220 0 net32
rlabel metal1 6670 10676 6670 10676 0 net33
rlabel metal1 8878 4658 8878 4658 0 net34
rlabel metal2 8970 7412 8970 7412 0 net35
rlabel metal1 5290 4012 5290 4012 0 net36
rlabel metal1 4738 3672 4738 3672 0 net37
rlabel metal1 4922 5746 4922 5746 0 net38
rlabel metal1 9292 7514 9292 7514 0 net39
rlabel metal1 8050 10676 8050 10676 0 net4
rlabel metal2 9246 6698 9246 6698 0 net40
rlabel metal1 8142 4658 8142 4658 0 net41
rlabel metal2 8326 4012 8326 4012 0 net42
rlabel via1 5098 10778 5098 10778 0 net5
rlabel metal1 3128 7854 3128 7854 0 net6
rlabel metal2 3450 5916 3450 5916 0 net7
rlabel metal1 4600 2618 4600 2618 0 net8
rlabel metal1 9936 2618 9936 2618 0 net9
rlabel metal2 6486 1588 6486 1588 0 op[0]
rlabel metal2 10442 7123 10442 7123 0 op[1]
rlabel metal2 10442 6239 10442 6239 0 op[2]
rlabel metal2 7774 959 7774 959 0 result[0]
rlabel metal2 7130 1520 7130 1520 0 result[1]
rlabel metal1 10580 8330 10580 8330 0 result[2]
rlabel metal1 6210 11322 6210 11322 0 result[3]
rlabel metal3 751 10268 751 10268 0 result[4]
rlabel metal3 1096 8228 1096 8228 0 result[5]
rlabel metal1 1426 5338 1426 5338 0 result[6]
rlabel metal3 751 3468 751 3468 0 result[7]
<< properties >>
string FIXED_BBOX 0 0 11998 14142
<< end >>
