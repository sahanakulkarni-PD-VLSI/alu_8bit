VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu_8bit
  CLASS BLOCK ;
  FOREIGN alu_8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 51.005 BY 61.725 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.965 10.640 14.565 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 22.855 10.640 24.455 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.745 10.640 34.345 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.635 10.640 44.235 49.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.140 45.320 19.740 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.660 45.320 29.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 37.180 45.320 38.780 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 46.700 45.320 48.300 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.665 10.640 11.265 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.555 10.640 21.155 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.445 10.640 31.045 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.335 10.640 40.935 49.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.840 45.320 16.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 24.360 45.320 25.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 33.880 45.320 35.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.400 45.320 45.000 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 10.240 51.005 10.840 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 20.440 51.005 21.040 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 40.840 51.005 41.440 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 57.725 29.350 61.725 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 17.040 51.005 17.640 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 23.840 51.005 24.440 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 44.240 51.005 44.840 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 57.725 26.130 61.725 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END b[7]
  PIN cin
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 13.640 51.005 14.240 ;
    END
  END cin
  PIN cout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END cout
  PIN op[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END op[0]
  PIN op[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 47.005 30.640 51.005 31.240 ;
    END
  END op[1]
  PIN op[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 47.005 34.040 51.005 34.640 ;
    END
  END op[2]
  PIN result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END result[0]
  PIN result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 27.240 51.005 27.840 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 47.005 37.440 51.005 38.040 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 57.725 22.910 61.725 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END result[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 45.270 49.045 ;
      LAYER li1 ;
        RECT 5.520 10.795 45.080 49.045 ;
      LAYER met1 ;
        RECT 4.210 9.560 45.930 49.200 ;
      LAYER met2 ;
        RECT 4.230 57.445 22.350 57.725 ;
        RECT 23.190 57.445 25.570 57.725 ;
        RECT 26.410 57.445 28.790 57.725 ;
        RECT 29.630 57.445 45.910 57.725 ;
        RECT 4.230 4.280 45.910 57.445 ;
        RECT 4.230 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 32.010 4.280 ;
        RECT 32.850 4.000 45.910 4.280 ;
      LAYER met3 ;
        RECT 3.750 48.640 47.005 49.125 ;
        RECT 4.400 47.240 47.005 48.640 ;
        RECT 3.750 45.240 47.005 47.240 ;
        RECT 4.400 43.840 46.605 45.240 ;
        RECT 3.750 41.840 47.005 43.840 ;
        RECT 4.400 40.440 46.605 41.840 ;
        RECT 3.750 38.440 47.005 40.440 ;
        RECT 4.400 37.040 46.605 38.440 ;
        RECT 3.750 35.040 47.005 37.040 ;
        RECT 4.400 33.640 46.605 35.040 ;
        RECT 3.750 31.640 47.005 33.640 ;
        RECT 4.400 30.240 46.605 31.640 ;
        RECT 3.750 28.240 47.005 30.240 ;
        RECT 4.400 26.840 46.605 28.240 ;
        RECT 3.750 24.840 47.005 26.840 ;
        RECT 4.400 23.440 46.605 24.840 ;
        RECT 3.750 21.440 47.005 23.440 ;
        RECT 3.750 20.040 46.605 21.440 ;
        RECT 3.750 18.040 47.005 20.040 ;
        RECT 4.400 16.640 46.605 18.040 ;
        RECT 3.750 14.640 47.005 16.640 ;
        RECT 3.750 13.240 46.605 14.640 ;
        RECT 3.750 11.240 47.005 13.240 ;
        RECT 3.750 9.840 46.605 11.240 ;
        RECT 3.750 9.695 47.005 9.840 ;
      LAYER met4 ;
        RECT 3.975 29.415 4.305 34.505 ;
  END
END alu_8bit
END LIBRARY

