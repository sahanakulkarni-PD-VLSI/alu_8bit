magic
tech sky130A
magscale 1 2
timestamp 1746634689
<< viali >>
rect 3407 10761 3441 10795
rect 4629 10761 4663 10795
rect 6561 10761 6595 10795
rect 3617 10693 3651 10727
rect 3801 10625 3835 10659
rect 3893 10625 3927 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4445 10625 4479 10659
rect 6009 10625 6043 10659
rect 6469 10625 6503 10659
rect 6929 10625 6963 10659
rect 8493 10625 8527 10659
rect 8677 10625 8711 10659
rect 9137 10625 9171 10659
rect 9413 10625 9447 10659
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 8217 10557 8251 10591
rect 3249 10489 3283 10523
rect 4813 10489 4847 10523
rect 7757 10489 7791 10523
rect 9045 10489 9079 10523
rect 9229 10489 9263 10523
rect 3433 10421 3467 10455
rect 4353 10421 4387 10455
rect 5825 10421 5859 10455
rect 6193 10421 6227 10455
rect 7113 10421 7147 10455
rect 8309 10421 8343 10455
rect 9137 10217 9171 10251
rect 3617 10081 3651 10115
rect 4629 10081 4663 10115
rect 5089 10081 5123 10115
rect 6193 10081 6227 10115
rect 6745 10081 6779 10115
rect 7573 10081 7607 10115
rect 8033 10081 8067 10115
rect 1409 10013 1443 10047
rect 4905 10013 4939 10047
rect 5549 10013 5583 10047
rect 5825 10013 5859 10047
rect 6561 10013 6595 10047
rect 7757 10013 7791 10047
rect 8125 10013 8159 10047
rect 8493 10013 8527 10047
rect 8677 10013 8711 10047
rect 8953 10013 8987 10047
rect 7113 9945 7147 9979
rect 1593 9877 1627 9911
rect 3157 9877 3191 9911
rect 6285 9877 6319 9911
rect 8585 9877 8619 9911
rect 3525 9673 3559 9707
rect 7665 9673 7699 9707
rect 8401 9673 8435 9707
rect 4873 9605 4907 9639
rect 5089 9605 5123 9639
rect 5733 9605 5767 9639
rect 7941 9605 7975 9639
rect 8151 9605 8185 9639
rect 2605 9537 2639 9571
rect 2789 9537 2823 9571
rect 3157 9537 3191 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 3801 9537 3835 9571
rect 3893 9537 3927 9571
rect 4629 9537 4663 9571
rect 5365 9537 5399 9571
rect 6009 9537 6043 9571
rect 6193 9537 6227 9571
rect 6561 9537 6595 9571
rect 6929 9537 6963 9571
rect 7021 9537 7055 9571
rect 7205 9537 7239 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 8309 9537 8343 9571
rect 8677 9537 8711 9571
rect 9045 9537 9079 9571
rect 9229 9537 9263 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 2881 9469 2915 9503
rect 5549 9469 5583 9503
rect 6377 9469 6411 9503
rect 7113 9469 7147 9503
rect 8585 9469 8619 9503
rect 8769 9469 8803 9503
rect 8861 9469 8895 9503
rect 9137 9469 9171 9503
rect 4169 9401 4203 9435
rect 5365 9401 5399 9435
rect 6837 9401 6871 9435
rect 2421 9333 2455 9367
rect 2789 9333 2823 9367
rect 2973 9333 3007 9367
rect 3065 9333 3099 9367
rect 3341 9333 3375 9367
rect 4721 9333 4755 9367
rect 4905 9333 4939 9367
rect 5825 9333 5859 9367
rect 9413 9333 9447 9367
rect 4445 9129 4479 9163
rect 1501 9061 1535 9095
rect 3525 9061 3559 9095
rect 9229 9061 9263 9095
rect 5365 8993 5399 9027
rect 8217 8993 8251 9027
rect 8309 8993 8343 9027
rect 1685 8925 1719 8959
rect 1777 8925 1811 8959
rect 2053 8925 2087 8959
rect 2145 8925 2179 8959
rect 2237 8925 2271 8959
rect 2421 8925 2455 8959
rect 2697 8925 2731 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 3801 8925 3835 8959
rect 4629 8925 4663 8959
rect 4905 8925 4939 8959
rect 5641 8925 5675 8959
rect 8401 8925 8435 8959
rect 8493 8925 8527 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9413 8925 9447 8959
rect 1935 8857 1969 8891
rect 3985 8857 4019 8891
rect 2513 8789 2547 8823
rect 4169 8789 4203 8823
rect 4813 8789 4847 8823
rect 8033 8789 8067 8823
rect 9045 8789 9079 8823
rect 1777 8585 1811 8619
rect 2237 8585 2271 8619
rect 5089 8517 5123 8551
rect 7573 8517 7607 8551
rect 7757 8517 7791 8551
rect 8861 8517 8895 8551
rect 1961 8449 1995 8483
rect 2145 8449 2179 8483
rect 2421 8449 2455 8483
rect 2513 8449 2547 8483
rect 2881 8449 2915 8483
rect 3801 8449 3835 8483
rect 4353 8449 4387 8483
rect 5273 8449 5307 8483
rect 5457 8449 5491 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 6929 8449 6963 8483
rect 7113 8449 7147 8483
rect 7481 8449 7515 8483
rect 7855 8449 7889 8483
rect 8033 8449 8067 8483
rect 8125 8449 8159 8483
rect 8217 8449 8251 8483
rect 9413 8449 9447 8483
rect 2789 8381 2823 8415
rect 3985 8381 4019 8415
rect 4261 8381 4295 8415
rect 7297 8313 7331 8347
rect 8493 8313 8527 8347
rect 5549 8245 5583 8279
rect 6377 8245 6411 8279
rect 7757 8245 7791 8279
rect 4813 8041 4847 8075
rect 7941 8041 7975 8075
rect 8493 8041 8527 8075
rect 6653 7973 6687 8007
rect 7665 7973 7699 8007
rect 7849 7905 7883 7939
rect 1409 7837 1443 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 5181 7837 5215 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 6101 7837 6135 7871
rect 6377 7837 6411 7871
rect 6469 7837 6503 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 7481 7837 7515 7871
rect 7757 7837 7791 7871
rect 8368 7837 8402 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 5273 7769 5307 7803
rect 6285 7769 6319 7803
rect 8244 7769 8278 7803
rect 1593 7701 1627 7735
rect 5089 7701 5123 7735
rect 5825 7701 5859 7735
rect 8677 7701 8711 7735
rect 9413 7701 9447 7735
rect 1777 7497 1811 7531
rect 3275 7497 3309 7531
rect 4277 7497 4311 7531
rect 4997 7497 5031 7531
rect 2329 7429 2363 7463
rect 3065 7429 3099 7463
rect 4077 7429 4111 7463
rect 5503 7429 5537 7463
rect 6653 7429 6687 7463
rect 7389 7429 7423 7463
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 2513 7361 2547 7395
rect 3525 7361 3559 7395
rect 3617 7361 3651 7395
rect 3801 7361 3835 7395
rect 5181 7361 5215 7395
rect 5273 7361 5307 7395
rect 5365 7361 5399 7395
rect 5641 7361 5675 7395
rect 7573 7361 7607 7395
rect 8861 7361 8895 7395
rect 9413 7361 9447 7395
rect 3985 7293 4019 7327
rect 7941 7293 7975 7327
rect 8125 7293 8159 7327
rect 3433 7225 3467 7259
rect 7021 7225 7055 7259
rect 1501 7157 1535 7191
rect 2145 7157 2179 7191
rect 3249 7157 3283 7191
rect 4261 7157 4295 7191
rect 4445 7157 4479 7191
rect 7113 7157 7147 7191
rect 8585 7157 8619 7191
rect 3893 6953 3927 6987
rect 4997 6953 5031 6987
rect 8677 6953 8711 6987
rect 8953 6817 8987 6851
rect 9137 6817 9171 6851
rect 9229 6817 9263 6851
rect 9321 6817 9355 6851
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 2329 6749 2363 6783
rect 2605 6749 2639 6783
rect 2789 6749 2823 6783
rect 2973 6749 3007 6783
rect 3249 6749 3283 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 4629 6749 4663 6783
rect 5457 6749 5491 6783
rect 7573 6749 7607 6783
rect 8217 6749 8251 6783
rect 8493 6749 8527 6783
rect 8769 6749 8803 6783
rect 9413 6749 9447 6783
rect 1777 6681 1811 6715
rect 2697 6681 2731 6715
rect 3433 6681 3467 6715
rect 1593 6613 1627 6647
rect 2053 6613 2087 6647
rect 2789 6613 2823 6647
rect 3065 6613 3099 6647
rect 4169 6613 4203 6647
rect 7389 6613 7423 6647
rect 7757 6613 7791 6647
rect 2329 6409 2363 6443
rect 7205 6409 7239 6443
rect 1843 6341 1877 6375
rect 2053 6341 2087 6375
rect 1409 6273 1443 6307
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2145 6273 2179 6307
rect 3341 6273 3375 6307
rect 3617 6273 3651 6307
rect 4169 6273 4203 6307
rect 4997 6273 5031 6307
rect 5549 6273 5583 6307
rect 5917 6273 5951 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 8401 6273 8435 6307
rect 8953 6273 8987 6307
rect 3801 6205 3835 6239
rect 4077 6205 4111 6239
rect 6377 6205 6411 6239
rect 8217 6205 8251 6239
rect 9229 6205 9263 6239
rect 1593 6137 1627 6171
rect 6837 6137 6871 6171
rect 7481 6137 7515 6171
rect 8493 6137 8527 6171
rect 3433 6069 3467 6103
rect 5089 6069 5123 6103
rect 6009 6069 6043 6103
rect 7757 6069 7791 6103
rect 1593 5865 1627 5899
rect 6101 5865 6135 5899
rect 9321 5865 9355 5899
rect 6193 5797 6227 5831
rect 8033 5797 8067 5831
rect 5457 5729 5491 5763
rect 6929 5729 6963 5763
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 4445 5661 4479 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 6377 5661 6411 5695
rect 6469 5661 6503 5695
rect 7113 5661 7147 5695
rect 7757 5661 7791 5695
rect 7895 5661 7929 5695
rect 8125 5661 8159 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 5615 5593 5649 5627
rect 5825 5593 5859 5627
rect 6745 5593 6779 5627
rect 6837 5593 6871 5627
rect 7297 5593 7331 5627
rect 9137 5593 9171 5627
rect 1685 5525 1719 5559
rect 4261 5525 4295 5559
rect 8309 5525 8343 5559
rect 1409 5321 1443 5355
rect 2145 5321 2179 5355
rect 3801 5321 3835 5355
rect 5457 5321 5491 5355
rect 6377 5321 6411 5355
rect 7297 5321 7331 5355
rect 1777 5253 1811 5287
rect 1915 5253 1949 5287
rect 2697 5253 2731 5287
rect 2789 5253 2823 5287
rect 3157 5253 3191 5287
rect 3357 5253 3391 5287
rect 5273 5253 5307 5287
rect 1593 5185 1627 5219
rect 1685 5185 1719 5219
rect 2421 5185 2455 5219
rect 4261 5185 4295 5219
rect 4445 5185 4479 5219
rect 4997 5185 5031 5219
rect 5733 5185 5767 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 7205 5185 7239 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 8401 5185 8435 5219
rect 8953 5185 8987 5219
rect 2053 5117 2087 5151
rect 2329 5117 2363 5151
rect 4905 5117 4939 5151
rect 5365 5117 5399 5151
rect 5641 5117 5675 5151
rect 5825 5117 5859 5151
rect 5917 5117 5951 5151
rect 4629 5049 4663 5083
rect 7021 5049 7055 5083
rect 8217 5049 8251 5083
rect 3341 4981 3375 5015
rect 3525 4981 3559 5015
rect 4077 4981 4111 5015
rect 4721 4981 4755 5015
rect 1501 4777 1535 4811
rect 1777 4777 1811 4811
rect 2881 4777 2915 4811
rect 5181 4777 5215 4811
rect 6745 4709 6779 4743
rect 7481 4709 7515 4743
rect 8493 4709 8527 4743
rect 4261 4641 4295 4675
rect 4721 4641 4755 4675
rect 1685 4573 1719 4607
rect 3249 4573 3283 4607
rect 3341 4573 3375 4607
rect 3525 4573 3559 4607
rect 3801 4573 3835 4607
rect 4353 4573 4387 4607
rect 4813 4573 4847 4607
rect 4997 4573 5031 4607
rect 6561 4573 6595 4607
rect 6837 4573 6871 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 8217 4573 8251 4607
rect 8493 4573 8527 4607
rect 9137 4573 9171 4607
rect 1961 4505 1995 4539
rect 2145 4505 2179 4539
rect 3065 4505 3099 4539
rect 7113 4505 7147 4539
rect 8953 4505 8987 4539
rect 9505 4505 9539 4539
rect 3433 4437 3467 4471
rect 3985 4437 4019 4471
rect 6929 4437 6963 4471
rect 6745 4233 6779 4267
rect 1409 4097 1443 4131
rect 4629 4097 4663 4131
rect 4997 4097 5031 4131
rect 5181 4097 5215 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 8585 4097 8619 4131
rect 9413 4097 9447 4131
rect 4905 4029 4939 4063
rect 6837 4029 6871 4063
rect 6929 4029 6963 4063
rect 7849 4029 7883 4063
rect 7941 4029 7975 4063
rect 8033 4029 8067 4063
rect 8125 4029 8159 4063
rect 8309 4029 8343 4063
rect 4813 3961 4847 3995
rect 7481 3961 7515 3995
rect 1593 3893 1627 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 6377 3893 6411 3927
rect 7665 3893 7699 3927
rect 9229 3893 9263 3927
rect 1869 3689 1903 3723
rect 2513 3689 2547 3723
rect 2789 3689 2823 3723
rect 3617 3689 3651 3723
rect 4721 3689 4755 3723
rect 5365 3689 5399 3723
rect 5917 3689 5951 3723
rect 6653 3689 6687 3723
rect 1961 3621 1995 3655
rect 2605 3621 2639 3655
rect 4905 3621 4939 3655
rect 9045 3621 9079 3655
rect 1777 3553 1811 3587
rect 2421 3553 2455 3587
rect 5825 3553 5859 3587
rect 8493 3553 8527 3587
rect 9505 3553 9539 3587
rect 2053 3485 2087 3519
rect 2513 3485 2547 3519
rect 3065 3485 3099 3519
rect 3157 3485 3191 3519
rect 3341 3485 3375 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4261 3485 4295 3519
rect 4997 3485 5031 3519
rect 5549 3485 5583 3519
rect 6929 3485 6963 3519
rect 7113 3485 7147 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 7941 3485 7975 3519
rect 8194 3485 8228 3519
rect 2973 3417 3007 3451
rect 4537 3417 4571 3451
rect 4753 3417 4787 3451
rect 5181 3417 5215 3451
rect 2145 3349 2179 3383
rect 2763 3349 2797 3383
rect 4169 3349 4203 3383
rect 6101 3349 6135 3383
rect 6837 3349 6871 3383
rect 3249 3145 3283 3179
rect 4261 3145 4295 3179
rect 4905 3145 4939 3179
rect 7021 3145 7055 3179
rect 7573 3145 7607 3179
rect 7849 3145 7883 3179
rect 9137 3145 9171 3179
rect 2881 3077 2915 3111
rect 4537 3077 4571 3111
rect 5733 3077 5767 3111
rect 8769 3077 8803 3111
rect 9045 3077 9079 3111
rect 4767 3043 4801 3077
rect 2697 3009 2731 3043
rect 2973 3009 3007 3043
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 4445 3009 4479 3043
rect 4997 3009 5031 3043
rect 5273 3009 5307 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 6653 3009 6687 3043
rect 7205 3009 7239 3043
rect 7573 3009 7607 3043
rect 7757 3009 7791 3043
rect 8401 3009 8435 3043
rect 8585 3009 8619 3043
rect 8953 3009 8987 3043
rect 5089 2941 5123 2975
rect 6101 2941 6135 2975
rect 6561 2941 6595 2975
rect 8309 2941 8343 2975
rect 9413 2941 9447 2975
rect 2697 2873 2731 2907
rect 7941 2873 7975 2907
rect 4445 2805 4479 2839
rect 4721 2805 4755 2839
rect 6377 2805 6411 2839
rect 3525 2601 3559 2635
rect 4169 2601 4203 2635
rect 5457 2601 5491 2635
rect 7941 2601 7975 2635
rect 8309 2601 8343 2635
rect 8677 2601 8711 2635
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5641 2397 5675 2431
rect 6469 2397 6503 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 7849 2397 7883 2431
rect 8033 2397 8067 2431
rect 8125 2397 8159 2431
rect 8493 2397 8527 2431
rect 5089 2329 5123 2363
rect 6837 2329 6871 2363
rect 7297 2261 7331 2295
rect 7573 2261 7607 2295
<< metal1 >>
rect 1104 10906 9844 10928
rect 1104 10854 2702 10906
rect 2754 10854 2766 10906
rect 2818 10854 2830 10906
rect 2882 10854 2894 10906
rect 2946 10854 2958 10906
rect 3010 10854 4887 10906
rect 4939 10854 4951 10906
rect 5003 10854 5015 10906
rect 5067 10854 5079 10906
rect 5131 10854 5143 10906
rect 5195 10854 7072 10906
rect 7124 10854 7136 10906
rect 7188 10854 7200 10906
rect 7252 10854 7264 10906
rect 7316 10854 7328 10906
rect 7380 10854 9257 10906
rect 9309 10854 9321 10906
rect 9373 10854 9385 10906
rect 9437 10854 9449 10906
rect 9501 10854 9513 10906
rect 9565 10854 9844 10906
rect 1104 10832 9844 10854
rect 3418 10801 3424 10804
rect 3395 10795 3424 10801
rect 3395 10761 3407 10795
rect 3476 10792 3482 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 3476 10764 4629 10792
rect 3395 10755 3424 10761
rect 3418 10752 3424 10755
rect 3476 10752 3482 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 4617 10755 4675 10761
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 5316 10764 6561 10792
rect 5316 10752 5322 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 6549 10755 6607 10761
rect 3605 10727 3663 10733
rect 3605 10693 3617 10727
rect 3651 10724 3663 10727
rect 3694 10724 3700 10736
rect 3651 10696 3700 10724
rect 3651 10693 3663 10696
rect 3605 10687 3663 10693
rect 3694 10684 3700 10696
rect 3752 10684 3758 10736
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4028 10696 4476 10724
rect 4028 10684 4034 10696
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3252 10628 3801 10656
rect 3252 10529 3280 10628
rect 3620 10600 3648 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 3602 10548 3608 10600
rect 3660 10548 3666 10600
rect 3896 10588 3924 10619
rect 4062 10616 4068 10668
rect 4120 10616 4126 10668
rect 4448 10665 4476 10696
rect 7742 10684 7748 10736
rect 7800 10724 7806 10736
rect 7800 10696 9444 10724
rect 7800 10684 7806 10696
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4172 10588 4200 10619
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5868 10628 6009 10656
rect 5868 10616 5874 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6457 10659 6515 10665
rect 6457 10656 6469 10659
rect 6144 10628 6469 10656
rect 6144 10616 6150 10628
rect 6457 10625 6469 10628
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6604 10628 6929 10656
rect 6604 10616 6610 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 8478 10616 8484 10668
rect 8536 10656 8542 10668
rect 8665 10659 8723 10665
rect 8536 10628 8616 10656
rect 8536 10616 8542 10628
rect 4614 10588 4620 10600
rect 3896 10560 4108 10588
rect 4172 10560 4620 10588
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10489 3295 10523
rect 4080 10520 4108 10560
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 5258 10548 5264 10600
rect 5316 10548 5322 10600
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7984 10560 8217 10588
rect 7984 10548 7990 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8588 10588 8616 10628
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 9122 10656 9128 10668
rect 8711 10628 9128 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 9416 10665 9444 10696
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 8588 10560 9260 10588
rect 8205 10551 8263 10557
rect 4801 10523 4859 10529
rect 4801 10520 4813 10523
rect 4080 10492 4813 10520
rect 3237 10483 3295 10489
rect 4801 10489 4813 10492
rect 4847 10489 4859 10523
rect 4801 10483 4859 10489
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7745 10523 7803 10529
rect 7745 10520 7757 10523
rect 6972 10492 7757 10520
rect 6972 10480 6978 10492
rect 7745 10489 7757 10492
rect 7791 10489 7803 10523
rect 7745 10483 7803 10489
rect 8110 10480 8116 10532
rect 8168 10520 8174 10532
rect 9232 10529 9260 10560
rect 9033 10523 9091 10529
rect 9033 10520 9045 10523
rect 8168 10492 9045 10520
rect 8168 10480 8174 10492
rect 9033 10489 9045 10492
rect 9079 10489 9091 10523
rect 9033 10483 9091 10489
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10489 9275 10523
rect 9217 10483 9275 10489
rect 3418 10412 3424 10464
rect 3476 10412 3482 10464
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4028 10424 4353 10452
rect 4028 10412 4034 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 5810 10412 5816 10464
rect 5868 10412 5874 10464
rect 6178 10412 6184 10464
rect 6236 10412 6242 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 7064 10424 7113 10452
rect 7064 10412 7070 10424
rect 7101 10421 7113 10424
rect 7147 10421 7159 10455
rect 7101 10415 7159 10421
rect 8294 10412 8300 10464
rect 8352 10412 8358 10464
rect 1104 10362 9844 10384
rect 1104 10310 2042 10362
rect 2094 10310 2106 10362
rect 2158 10310 2170 10362
rect 2222 10310 2234 10362
rect 2286 10310 2298 10362
rect 2350 10310 4227 10362
rect 4279 10310 4291 10362
rect 4343 10310 4355 10362
rect 4407 10310 4419 10362
rect 4471 10310 4483 10362
rect 4535 10310 6412 10362
rect 6464 10310 6476 10362
rect 6528 10310 6540 10362
rect 6592 10310 6604 10362
rect 6656 10310 6668 10362
rect 6720 10310 8597 10362
rect 8649 10310 8661 10362
rect 8713 10310 8725 10362
rect 8777 10310 8789 10362
rect 8841 10310 8853 10362
rect 8905 10310 9844 10362
rect 1104 10288 9844 10310
rect 9122 10208 9128 10260
rect 9180 10208 9186 10260
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 5316 10152 7604 10180
rect 5316 10140 5322 10152
rect 3602 10072 3608 10124
rect 3660 10072 3666 10124
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4522 10112 4528 10124
rect 3752 10084 4528 10112
rect 3752 10072 3758 10084
rect 4522 10072 4528 10084
rect 4580 10112 4586 10124
rect 4617 10115 4675 10121
rect 4617 10112 4629 10115
rect 4580 10084 4629 10112
rect 4580 10072 4586 10084
rect 4617 10081 4629 10084
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5350 10112 5356 10124
rect 5123 10084 5356 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 6196 10121 6224 10152
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 7576 10121 7604 10152
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7984 10084 8033 10112
rect 7984 10072 7990 10084
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8444 10084 8984 10112
rect 8444 10072 8450 10084
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4154 10044 4160 10056
rect 4028 10016 4160 10044
rect 4028 10004 4034 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4856 10016 4905 10044
rect 4856 10004 4862 10016
rect 4893 10013 4905 10016
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 5994 10044 6000 10056
rect 5859 10016 6000 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 5552 9976 5580 10007
rect 5994 10004 6000 10016
rect 6052 10044 6058 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6052 10016 6561 10044
rect 6052 10004 6058 10016
rect 6549 10013 6561 10016
rect 6595 10044 6607 10047
rect 7006 10044 7012 10056
rect 6595 10016 7012 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7006 10004 7012 10016
rect 7064 10044 7070 10056
rect 7466 10044 7472 10056
rect 7064 10016 7472 10044
rect 7064 10004 7070 10016
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 6730 9976 6736 9988
rect 5552 9948 6736 9976
rect 6730 9936 6736 9948
rect 6788 9976 6794 9988
rect 7101 9979 7159 9985
rect 7101 9976 7113 9979
rect 6788 9948 7113 9976
rect 6788 9936 6794 9948
rect 7101 9945 7113 9948
rect 7147 9945 7159 9979
rect 8128 9976 8156 10007
rect 8478 10004 8484 10056
rect 8536 10004 8542 10056
rect 8956 10053 8984 10084
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 8386 9976 8392 9988
rect 8128 9948 8392 9976
rect 7101 9939 7159 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 8680 9976 8708 10007
rect 9122 9976 9128 9988
rect 8680 9948 9128 9976
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 2590 9908 2596 9920
rect 1627 9880 2596 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 6270 9868 6276 9920
rect 6328 9868 6334 9920
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 8662 9908 8668 9920
rect 8619 9880 8668 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 1104 9818 9844 9840
rect 1104 9766 2702 9818
rect 2754 9766 2766 9818
rect 2818 9766 2830 9818
rect 2882 9766 2894 9818
rect 2946 9766 2958 9818
rect 3010 9766 4887 9818
rect 4939 9766 4951 9818
rect 5003 9766 5015 9818
rect 5067 9766 5079 9818
rect 5131 9766 5143 9818
rect 5195 9766 7072 9818
rect 7124 9766 7136 9818
rect 7188 9766 7200 9818
rect 7252 9766 7264 9818
rect 7316 9766 7328 9818
rect 7380 9766 9257 9818
rect 9309 9766 9321 9818
rect 9373 9766 9385 9818
rect 9437 9766 9449 9818
rect 9501 9766 9513 9818
rect 9565 9766 9844 9818
rect 1104 9744 9844 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3513 9707 3571 9713
rect 3513 9704 3525 9707
rect 3476 9676 3525 9704
rect 3476 9664 3482 9676
rect 3513 9673 3525 9676
rect 3559 9704 3571 9707
rect 7653 9707 7711 9713
rect 3559 9676 3924 9704
rect 3559 9673 3571 9676
rect 3513 9667 3571 9673
rect 3896 9636 3924 9676
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 7742 9704 7748 9716
rect 7699 9676 7748 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 8386 9664 8392 9716
rect 8444 9664 8450 9716
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 8536 9676 9260 9704
rect 8536 9664 8542 9676
rect 2608 9608 3832 9636
rect 3896 9608 4752 9636
rect 2608 9580 2636 9608
rect 2590 9528 2596 9580
rect 2648 9528 2654 9580
rect 2774 9528 2780 9580
rect 2832 9528 2838 9580
rect 2884 9509 2912 9608
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3804 9577 3832 9608
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4062 9568 4068 9580
rect 3927 9540 4068 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9469 2927 9503
rect 2869 9463 2927 9469
rect 3160 9432 3188 9528
rect 3620 9500 3648 9531
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4580 9540 4629 9568
rect 4580 9528 4586 9540
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4724 9568 4752 9608
rect 4798 9596 4804 9648
rect 4856 9645 4862 9648
rect 4856 9639 4919 9645
rect 4856 9605 4873 9639
rect 4907 9605 4919 9639
rect 4856 9599 4919 9605
rect 5077 9639 5135 9645
rect 5077 9605 5089 9639
rect 5123 9605 5135 9639
rect 5077 9599 5135 9605
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 6270 9636 6276 9648
rect 5767 9608 6276 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 4856 9596 4862 9599
rect 5092 9568 5120 9599
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 7929 9639 7987 9645
rect 7929 9636 7941 9639
rect 6380 9608 7052 9636
rect 4724 9540 5120 9568
rect 4617 9531 4675 9537
rect 3620 9472 4200 9500
rect 4172 9441 4200 9472
rect 5092 9444 5120 9540
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6380 9568 6408 9608
rect 6236 9540 6408 9568
rect 6549 9571 6607 9577
rect 6236 9528 6242 9540
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 6730 9568 6736 9580
rect 6595 9540 6736 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7024 9577 7052 9608
rect 7760 9608 7941 9636
rect 7760 9580 7788 9608
rect 7929 9605 7941 9608
rect 7975 9605 7987 9639
rect 7929 9599 7987 9605
rect 8110 9596 8116 9648
rect 8168 9645 8174 9648
rect 8168 9639 8197 9645
rect 8185 9605 8197 9639
rect 8168 9599 8197 9605
rect 8168 9596 8174 9599
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 7466 9568 7472 9580
rect 7239 9540 7472 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 7883 9540 7917 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 6196 9500 6224 9528
rect 5592 9472 6224 9500
rect 6365 9503 6423 9509
rect 5592 9460 5598 9472
rect 6365 9469 6377 9503
rect 6411 9500 6423 9503
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 6411 9472 7113 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 2792 9404 3188 9432
rect 4157 9435 4215 9441
rect 2406 9324 2412 9376
rect 2464 9324 2470 9376
rect 2792 9373 2820 9404
rect 4157 9401 4169 9435
rect 4203 9401 4215 9435
rect 4157 9395 4215 9401
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 5132 9404 5365 9432
rect 5132 9392 5138 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 6178 9392 6184 9444
rect 6236 9432 6242 9444
rect 6380 9432 6408 9463
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7852 9500 7880 9531
rect 8018 9528 8024 9580
rect 8076 9528 8082 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8496 9568 8524 9664
rect 9122 9596 9128 9648
rect 9180 9596 9186 9648
rect 8343 9540 8524 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9140 9568 9168 9596
rect 9232 9577 9260 9676
rect 9079 9540 9168 9568
rect 9217 9571 9275 9577
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 7708 9472 8585 9500
rect 7708 9460 7714 9472
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8895 9472 9137 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 6236 9404 6408 9432
rect 6236 9392 6242 9404
rect 6822 9392 6828 9444
rect 6880 9392 6886 9444
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 8018 9432 8024 9444
rect 7524 9404 8024 9432
rect 7524 9392 7530 9404
rect 8018 9392 8024 9404
rect 8076 9392 8082 9444
rect 8202 9392 8208 9444
rect 8260 9432 8266 9444
rect 9508 9432 9536 9531
rect 8260 9404 9536 9432
rect 8260 9392 8266 9404
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9333 2835 9367
rect 2777 9327 2835 9333
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3329 9367 3387 9373
rect 3329 9364 3341 9367
rect 3108 9336 3341 9364
rect 3108 9324 3114 9336
rect 3329 9333 3341 9336
rect 3375 9333 3387 9367
rect 3329 9327 3387 9333
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 4890 9324 4896 9376
rect 4948 9324 4954 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5813 9367 5871 9373
rect 5813 9364 5825 9367
rect 5500 9336 5825 9364
rect 5500 9324 5506 9336
rect 5813 9333 5825 9336
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8110 9364 8116 9376
rect 7800 9336 8116 9364
rect 7800 9324 7806 9336
rect 8110 9324 8116 9336
rect 8168 9364 8174 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 8168 9336 9413 9364
rect 8168 9324 8174 9336
rect 9401 9333 9413 9336
rect 9447 9364 9459 9367
rect 9582 9364 9588 9376
rect 9447 9336 9588 9364
rect 9447 9333 9459 9336
rect 9401 9327 9459 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 1104 9274 9844 9296
rect 1104 9222 2042 9274
rect 2094 9222 2106 9274
rect 2158 9222 2170 9274
rect 2222 9222 2234 9274
rect 2286 9222 2298 9274
rect 2350 9222 4227 9274
rect 4279 9222 4291 9274
rect 4343 9222 4355 9274
rect 4407 9222 4419 9274
rect 4471 9222 4483 9274
rect 4535 9222 6412 9274
rect 6464 9222 6476 9274
rect 6528 9222 6540 9274
rect 6592 9222 6604 9274
rect 6656 9222 6668 9274
rect 6720 9222 8597 9274
rect 8649 9222 8661 9274
rect 8713 9222 8725 9274
rect 8777 9222 8789 9274
rect 8841 9222 8853 9274
rect 8905 9222 9844 9274
rect 1104 9200 9844 9222
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4614 9160 4620 9172
rect 4479 9132 4620 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1489 9095 1547 9101
rect 1489 9092 1501 9095
rect 900 9064 1501 9092
rect 900 9052 906 9064
rect 1489 9061 1501 9064
rect 1535 9061 1547 9095
rect 1489 9055 1547 9061
rect 2406 9052 2412 9104
rect 2464 9052 2470 9104
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 3513 9095 3571 9101
rect 3513 9092 3525 9095
rect 2556 9064 3525 9092
rect 2556 9052 2562 9064
rect 3513 9061 3525 9064
rect 3559 9092 3571 9095
rect 4890 9092 4896 9104
rect 3559 9064 4896 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 9217 9095 9275 9101
rect 9217 9092 9229 9095
rect 7616 9064 9229 9092
rect 7616 9052 7622 9064
rect 9217 9061 9229 9064
rect 9263 9061 9275 9095
rect 9217 9055 9275 9061
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2424 9024 2452 9052
rect 1912 8996 2084 9024
rect 1912 8984 1918 8996
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1688 8820 1716 8919
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 2056 8965 2084 8996
rect 2148 8996 2452 9024
rect 2148 8965 2176 8996
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 5353 9027 5411 9033
rect 2648 8996 3832 9024
rect 2648 8984 2654 8996
rect 3436 8965 3464 8996
rect 3804 8965 3832 8996
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 5810 9024 5816 9036
rect 5399 8996 5816 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 8202 8984 8208 9036
rect 8260 8984 8266 9036
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8570 9024 8576 9036
rect 8343 8996 8576 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8956 2467 8959
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2455 8928 2697 8956
rect 2455 8925 2467 8928
rect 2409 8919 2467 8925
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 1946 8897 1952 8900
rect 1923 8891 1952 8897
rect 1923 8857 1935 8891
rect 1923 8851 1952 8857
rect 1946 8848 1952 8851
rect 2004 8848 2010 8900
rect 2240 8888 2268 8919
rect 2958 8888 2964 8900
rect 2240 8860 2964 8888
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 3326 8848 3332 8900
rect 3384 8888 3390 8900
rect 3620 8888 3648 8919
rect 3973 8891 4031 8897
rect 3973 8888 3985 8891
rect 3384 8860 3985 8888
rect 3384 8848 3390 8860
rect 3973 8857 3985 8860
rect 4019 8888 4031 8891
rect 4632 8888 4660 8919
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4856 8928 4905 8956
rect 4856 8916 4862 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8956 5687 8959
rect 5718 8956 5724 8968
rect 5675 8928 5724 8956
rect 5675 8925 5687 8928
rect 5629 8919 5687 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8312 8956 8340 8987
rect 8570 8984 8576 8996
rect 8628 9024 8634 9036
rect 9306 9024 9312 9036
rect 8628 8996 9312 9024
rect 8628 8984 8634 8996
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 7892 8928 8340 8956
rect 7892 8916 7898 8928
rect 8386 8916 8392 8968
rect 8444 8916 8450 8968
rect 8478 8916 8484 8968
rect 8536 8916 8542 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 9088 8928 9137 8956
rect 9088 8916 9094 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 9272 8928 9413 8956
rect 9272 8916 9278 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 4019 8860 4660 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 1688 8792 2513 8820
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 3844 8792 4169 8820
rect 3844 8780 3850 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4157 8783 4215 8789
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8820 4859 8823
rect 5074 8820 5080 8832
rect 4847 8792 5080 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8260 8792 9045 8820
rect 8260 8780 8266 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 9033 8783 9091 8789
rect 1104 8730 9844 8752
rect 1104 8678 2702 8730
rect 2754 8678 2766 8730
rect 2818 8678 2830 8730
rect 2882 8678 2894 8730
rect 2946 8678 2958 8730
rect 3010 8678 4887 8730
rect 4939 8678 4951 8730
rect 5003 8678 5015 8730
rect 5067 8678 5079 8730
rect 5131 8678 5143 8730
rect 5195 8678 7072 8730
rect 7124 8678 7136 8730
rect 7188 8678 7200 8730
rect 7252 8678 7264 8730
rect 7316 8678 7328 8730
rect 7380 8678 9257 8730
rect 9309 8678 9321 8730
rect 9373 8678 9385 8730
rect 9437 8678 9449 8730
rect 9501 8678 9513 8730
rect 9565 8678 9844 8730
rect 1104 8656 9844 8678
rect 1762 8576 1768 8628
rect 1820 8576 1826 8628
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 2004 8588 2237 8616
rect 2004 8576 2010 8588
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 2225 8579 2283 8585
rect 7466 8576 7472 8628
rect 7524 8576 7530 8628
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 8570 8616 8576 8628
rect 8220 8588 8576 8616
rect 2424 8520 3924 8548
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 2424 8489 2452 8520
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1360 8452 1961 8480
rect 1360 8440 1366 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2148 8412 2176 8443
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 3786 8480 3792 8492
rect 2915 8452 3792 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 2516 8412 2544 8440
rect 2148 8384 2544 8412
rect 2590 8372 2596 8424
rect 2648 8412 2654 8424
rect 2777 8415 2835 8421
rect 2777 8412 2789 8415
rect 2648 8384 2789 8412
rect 2648 8372 2654 8384
rect 2777 8381 2789 8384
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 3896 8344 3924 8520
rect 4798 8508 4804 8560
rect 4856 8548 4862 8560
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 4856 8520 5089 8548
rect 4856 8508 4862 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 6822 8548 6828 8560
rect 5077 8511 5135 8517
rect 5276 8520 6828 8548
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4706 8480 4712 8492
rect 4387 8452 4712 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5276 8489 5304 8520
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7484 8548 7512 8576
rect 7561 8551 7619 8557
rect 7561 8548 7573 8551
rect 7484 8520 7573 8548
rect 7561 8517 7573 8520
rect 7607 8517 7619 8551
rect 7561 8511 7619 8517
rect 7745 8551 7803 8557
rect 7745 8517 7757 8551
rect 7791 8548 7803 8551
rect 8128 8548 8156 8576
rect 7791 8520 8156 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4798 8412 4804 8424
rect 4295 8384 4804 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 5534 8412 5540 8424
rect 5132 8384 5540 8412
rect 5132 8372 5138 8384
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 5736 8412 5764 8443
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5868 8452 5917 8480
rect 5868 8440 5874 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6546 8480 6552 8492
rect 6328 8452 6552 8480
rect 6328 8440 6334 8452
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 5592 8384 5764 8412
rect 5592 8372 5598 8384
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 6748 8412 6776 8443
rect 6236 8384 6776 8412
rect 6236 8372 6242 8384
rect 5994 8344 6000 8356
rect 3896 8316 6000 8344
rect 5994 8304 6000 8316
rect 6052 8344 6058 8356
rect 6932 8344 6960 8443
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 7064 8452 7113 8480
rect 7064 8440 7070 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 7469 8483 7527 8489
rect 7843 8483 7901 8489
rect 7469 8480 7481 8483
rect 7432 8452 7481 8480
rect 7432 8440 7438 8452
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7668 8455 7855 8483
rect 7668 8412 7696 8455
rect 7843 8449 7855 8455
rect 7889 8449 7901 8483
rect 7843 8443 7901 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 7208 8384 7696 8412
rect 8036 8412 8064 8443
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 8220 8489 8248 8588
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 8294 8508 8300 8560
rect 8352 8508 8358 8560
rect 8386 8508 8392 8560
rect 8444 8548 8450 8560
rect 8849 8551 8907 8557
rect 8849 8548 8861 8551
rect 8444 8520 8861 8548
rect 8444 8508 8450 8520
rect 8849 8517 8861 8520
rect 8895 8517 8907 8551
rect 8849 8511 8907 8517
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8312 8412 8340 8508
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 8036 8384 8340 8412
rect 7098 8344 7104 8356
rect 6052 8316 7104 8344
rect 6052 8304 6058 8316
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5442 8276 5448 8288
rect 5224 8248 5448 8276
rect 5224 8236 5230 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5534 8236 5540 8288
rect 5592 8236 5598 8288
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 5684 8248 6377 8276
rect 5684 8236 5690 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6365 8239 6423 8245
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 7208 8276 7236 8384
rect 7285 8347 7343 8353
rect 7285 8313 7297 8347
rect 7331 8344 7343 8347
rect 8294 8344 8300 8356
rect 7331 8316 7512 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 6604 8248 7236 8276
rect 7484 8276 7512 8316
rect 7668 8316 8300 8344
rect 7668 8276 7696 8316
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 8478 8304 8484 8356
rect 8536 8304 8542 8356
rect 7484 8248 7696 8276
rect 7745 8279 7803 8285
rect 6604 8236 6610 8248
rect 7745 8245 7757 8279
rect 7791 8276 7803 8279
rect 9030 8276 9036 8288
rect 7791 8248 9036 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 1104 8186 9844 8208
rect 1104 8134 2042 8186
rect 2094 8134 2106 8186
rect 2158 8134 2170 8186
rect 2222 8134 2234 8186
rect 2286 8134 2298 8186
rect 2350 8134 4227 8186
rect 4279 8134 4291 8186
rect 4343 8134 4355 8186
rect 4407 8134 4419 8186
rect 4471 8134 4483 8186
rect 4535 8134 6412 8186
rect 6464 8134 6476 8186
rect 6528 8134 6540 8186
rect 6592 8134 6604 8186
rect 6656 8134 6668 8186
rect 6720 8134 8597 8186
rect 8649 8134 8661 8186
rect 8713 8134 8725 8186
rect 8777 8134 8789 8186
rect 8841 8134 8853 8186
rect 8905 8134 9844 8186
rect 1104 8112 9844 8134
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 6086 8072 6092 8084
rect 4847 8044 6092 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 7929 8075 7987 8081
rect 7929 8041 7941 8075
rect 7975 8072 7987 8075
rect 8018 8072 8024 8084
rect 7975 8044 8024 8072
rect 7975 8041 7987 8044
rect 7929 8035 7987 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 9122 8072 9128 8084
rect 8527 8044 9128 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 6641 8007 6699 8013
rect 6641 8004 6653 8007
rect 4816 7976 6653 8004
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 4614 7828 4620 7880
rect 4672 7828 4678 7880
rect 2590 7760 2596 7812
rect 2648 7800 2654 7812
rect 4816 7800 4844 7976
rect 6641 7973 6653 7976
rect 6687 7973 6699 8007
rect 6641 7967 6699 7973
rect 7653 8007 7711 8013
rect 7653 7973 7665 8007
rect 7699 8004 7711 8007
rect 8110 8004 8116 8016
rect 7699 7976 8116 8004
rect 7699 7973 7711 7976
rect 7653 7967 7711 7973
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8294 7964 8300 8016
rect 8352 7964 8358 8016
rect 5718 7936 5724 7948
rect 4908 7908 5724 7936
rect 4908 7877 4936 7908
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7837 7939 7895 7945
rect 6380 7908 7512 7936
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 5994 7868 6000 7880
rect 5675 7840 6000 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 2648 7772 5273 7800
rect 2648 7760 2654 7772
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 5552 7800 5580 7831
rect 5994 7828 6000 7840
rect 6052 7868 6058 7880
rect 6380 7877 6408 7908
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 6052 7840 6101 7868
rect 6052 7828 6058 7840
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6503 7840 6684 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6178 7800 6184 7812
rect 5552 7772 6184 7800
rect 5261 7763 5319 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6270 7760 6276 7812
rect 6328 7760 6334 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 3786 7732 3792 7744
rect 1627 7704 3792 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 5350 7732 5356 7744
rect 5123 7704 5356 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5810 7692 5816 7744
rect 5868 7692 5874 7744
rect 6656 7732 6684 7840
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7484 7877 7512 7908
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8202 7936 8208 7948
rect 7883 7908 8208 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8312 7936 8340 7964
rect 8312 7908 8616 7936
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7484 7800 7512 7831
rect 7742 7828 7748 7880
rect 7800 7828 7806 7880
rect 8386 7877 8392 7880
rect 8356 7871 8392 7877
rect 8356 7868 8368 7871
rect 7852 7840 8368 7868
rect 7852 7800 7880 7840
rect 8356 7837 8368 7840
rect 8356 7831 8392 7837
rect 8386 7828 8392 7831
rect 8444 7828 8450 7880
rect 8588 7877 8616 7908
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9030 7868 9036 7880
rect 8987 7840 9036 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 7484 7772 7880 7800
rect 8232 7803 8290 7809
rect 8232 7769 8244 7803
rect 8278 7800 8290 7803
rect 8588 7800 8616 7831
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 8278 7772 8616 7800
rect 8278 7769 8290 7772
rect 8232 7763 8290 7769
rect 8665 7735 8723 7741
rect 8665 7732 8677 7735
rect 6656 7704 8677 7732
rect 8665 7701 8677 7704
rect 8711 7701 8723 7735
rect 8665 7695 8723 7701
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9180 7704 9413 7732
rect 9180 7692 9186 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 1104 7642 9844 7664
rect 1104 7590 2702 7642
rect 2754 7590 2766 7642
rect 2818 7590 2830 7642
rect 2882 7590 2894 7642
rect 2946 7590 2958 7642
rect 3010 7590 4887 7642
rect 4939 7590 4951 7642
rect 5003 7590 5015 7642
rect 5067 7590 5079 7642
rect 5131 7590 5143 7642
rect 5195 7590 7072 7642
rect 7124 7590 7136 7642
rect 7188 7590 7200 7642
rect 7252 7590 7264 7642
rect 7316 7590 7328 7642
rect 7380 7590 9257 7642
rect 9309 7590 9321 7642
rect 9373 7590 9385 7642
rect 9437 7590 9449 7642
rect 9501 7590 9513 7642
rect 9565 7590 9844 7642
rect 1104 7568 9844 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7497 1823 7531
rect 1765 7491 1823 7497
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 1780 7392 1808 7491
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3263 7531 3321 7537
rect 3263 7528 3275 7531
rect 2740 7500 3275 7528
rect 2740 7488 2746 7500
rect 3263 7497 3275 7500
rect 3309 7528 3321 7531
rect 3878 7528 3884 7540
rect 3309 7500 3884 7528
rect 3309 7497 3321 7500
rect 3263 7491 3321 7497
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 3970 7488 3976 7540
rect 4028 7528 4034 7540
rect 4265 7531 4323 7537
rect 4265 7528 4277 7531
rect 4028 7500 4277 7528
rect 4028 7488 4034 7500
rect 4265 7497 4277 7500
rect 4311 7497 4323 7531
rect 4265 7491 4323 7497
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 4672 7500 4997 7528
rect 4672 7488 4678 7500
rect 4985 7497 4997 7500
rect 5031 7497 5043 7531
rect 4985 7491 5043 7497
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 2317 7463 2375 7469
rect 2317 7429 2329 7463
rect 2363 7460 2375 7463
rect 2406 7460 2412 7472
rect 2363 7432 2412 7460
rect 2363 7429 2375 7432
rect 2317 7423 2375 7429
rect 2406 7420 2412 7432
rect 2464 7420 2470 7472
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7429 3111 7463
rect 3988 7460 4016 7488
rect 3053 7423 3111 7429
rect 3528 7432 4016 7460
rect 4065 7463 4123 7469
rect 1719 7364 1808 7392
rect 1949 7395 2007 7401
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3068 7392 3096 7423
rect 3528 7401 3556 7432
rect 4065 7429 4077 7463
rect 4111 7429 4123 7463
rect 5368 7460 5396 7488
rect 4065 7423 4123 7429
rect 5184 7432 5396 7460
rect 5491 7463 5549 7469
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2547 7364 2774 7392
rect 3068 7364 3525 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 1964 7324 1992 7355
rect 2406 7324 2412 7336
rect 1964 7296 2412 7324
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2746 7324 2774 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3050 7324 3056 7336
rect 2746 7296 3056 7324
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 3620 7324 3648 7355
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 4080 7392 4108 7423
rect 5184 7401 5212 7432
rect 5491 7429 5503 7463
rect 5537 7460 5549 7463
rect 5810 7460 5816 7472
rect 5537 7432 5816 7460
rect 5537 7429 5549 7432
rect 5491 7423 5549 7429
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 7377 7463 7435 7469
rect 7377 7460 7389 7463
rect 6687 7432 7389 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 7377 7429 7389 7432
rect 7423 7460 7435 7463
rect 8386 7460 8392 7472
rect 7423 7432 8392 7460
rect 7423 7429 7435 7432
rect 7377 7423 7435 7429
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 3844 7364 4108 7392
rect 5169 7395 5227 7401
rect 3844 7352 3850 7364
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 3344 7296 3648 7324
rect 3973 7327 4031 7333
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 2004 7160 2145 7188
rect 2004 7148 2010 7160
rect 2133 7157 2145 7160
rect 2179 7157 2191 7191
rect 2133 7151 2191 7157
rect 3237 7191 3295 7197
rect 3237 7157 3249 7191
rect 3283 7188 3295 7191
rect 3344 7188 3372 7296
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4706 7324 4712 7336
rect 4019 7296 4712 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5276 7324 5304 7355
rect 5350 7352 5356 7404
rect 5408 7352 5414 7404
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 7607 7364 8861 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 8849 7361 8861 7364
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 5534 7324 5540 7336
rect 5276 7296 5540 7324
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 3421 7259 3479 7265
rect 3421 7225 3433 7259
rect 3467 7256 3479 7259
rect 4154 7256 4160 7268
rect 3467 7228 4160 7256
rect 3467 7225 3479 7228
rect 3421 7219 3479 7225
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 6972 7228 7021 7256
rect 6972 7216 6978 7228
rect 7009 7225 7021 7228
rect 7055 7256 7067 7259
rect 7576 7256 7604 7355
rect 9398 7352 9404 7404
rect 9456 7352 9462 7404
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8018 7324 8024 7336
rect 7975 7296 8024 7324
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8294 7324 8300 7336
rect 8159 7296 8300 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 7055 7228 7604 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 4246 7188 4252 7200
rect 3283 7160 4252 7188
rect 3283 7157 3295 7160
rect 3237 7151 3295 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4798 7188 4804 7200
rect 4479 7160 4804 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 7101 7191 7159 7197
rect 7101 7188 7113 7191
rect 6328 7160 7113 7188
rect 6328 7148 6334 7160
rect 7101 7157 7113 7160
rect 7147 7157 7159 7191
rect 7101 7151 7159 7157
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 8128 7188 8156 7287
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 7524 7160 8156 7188
rect 8573 7191 8631 7197
rect 7524 7148 7530 7160
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 9214 7188 9220 7200
rect 8619 7160 9220 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 1104 7098 9844 7120
rect 1104 7046 2042 7098
rect 2094 7046 2106 7098
rect 2158 7046 2170 7098
rect 2222 7046 2234 7098
rect 2286 7046 2298 7098
rect 2350 7046 4227 7098
rect 4279 7046 4291 7098
rect 4343 7046 4355 7098
rect 4407 7046 4419 7098
rect 4471 7046 4483 7098
rect 4535 7046 6412 7098
rect 6464 7046 6476 7098
rect 6528 7046 6540 7098
rect 6592 7046 6604 7098
rect 6656 7046 6668 7098
rect 6720 7046 8597 7098
rect 8649 7046 8661 7098
rect 8713 7046 8725 7098
rect 8777 7046 8789 7098
rect 8841 7046 8853 7098
rect 8905 7046 9844 7098
rect 1104 7024 9844 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 1912 6956 3832 6984
rect 1912 6944 1918 6956
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 2498 6916 2504 6928
rect 1636 6888 2504 6916
rect 1636 6876 1642 6888
rect 2498 6876 2504 6888
rect 2556 6916 2562 6928
rect 3804 6916 3832 6956
rect 3878 6944 3884 6996
rect 3936 6944 3942 6996
rect 4985 6987 5043 6993
rect 4985 6953 4997 6987
rect 5031 6984 5043 6987
rect 5442 6984 5448 6996
rect 5031 6956 5448 6984
rect 5031 6953 5043 6956
rect 4985 6947 5043 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 8665 6987 8723 6993
rect 8665 6953 8677 6987
rect 8711 6984 8723 6987
rect 9030 6984 9036 6996
rect 8711 6956 9036 6984
rect 8711 6953 8723 6956
rect 8665 6947 8723 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 5350 6916 5356 6928
rect 2556 6888 2820 6916
rect 3804 6888 5356 6916
rect 2556 6876 2562 6888
rect 2682 6848 2688 6860
rect 1964 6820 2688 6848
rect 1964 6789 1992 6820
rect 2332 6789 2360 6820
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 2792 6848 2820 6888
rect 5350 6876 5356 6888
rect 5408 6916 5414 6928
rect 5534 6916 5540 6928
rect 5408 6888 5540 6916
rect 5408 6876 5414 6888
rect 5534 6876 5540 6888
rect 5592 6916 5598 6928
rect 6730 6916 6736 6928
rect 5592 6888 6736 6916
rect 5592 6876 5598 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 2792 6820 3188 6848
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 1765 6715 1823 6721
rect 1765 6712 1777 6715
rect 1360 6684 1777 6712
rect 1360 6672 1366 6684
rect 1765 6681 1777 6684
rect 1811 6681 1823 6715
rect 2240 6712 2268 6743
rect 2590 6740 2596 6792
rect 2648 6740 2654 6792
rect 2792 6789 2820 6820
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6780 3019 6783
rect 3050 6780 3056 6792
rect 3007 6752 3056 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 2498 6712 2504 6724
rect 2240 6684 2504 6712
rect 1765 6675 1823 6681
rect 2498 6672 2504 6684
rect 2556 6672 2562 6724
rect 2685 6715 2743 6721
rect 2685 6681 2697 6715
rect 2731 6712 2743 6715
rect 3160 6712 3188 6820
rect 3252 6820 3924 6848
rect 3252 6789 3280 6820
rect 3896 6792 3924 6820
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 9122 6808 9128 6860
rect 9180 6808 9186 6860
rect 9214 6808 9220 6860
rect 9272 6808 9278 6860
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9582 6848 9588 6860
rect 9355 6820 9588 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3237 6743 3295 6749
rect 3436 6752 3801 6780
rect 3326 6712 3332 6724
rect 2731 6684 3096 6712
rect 3160 6684 3332 6712
rect 2731 6681 2743 6684
rect 2685 6675 2743 6681
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1670 6644 1676 6656
rect 1627 6616 1676 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2041 6647 2099 6653
rect 2041 6644 2053 6647
rect 1912 6616 2053 6644
rect 1912 6604 1918 6616
rect 2041 6613 2053 6616
rect 2087 6613 2099 6647
rect 2041 6607 2099 6613
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 3068 6653 3096 6684
rect 3326 6672 3332 6684
rect 3384 6712 3390 6724
rect 3436 6721 3464 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4304 6752 4629 6780
rect 4304 6740 4310 6752
rect 4617 6749 4629 6752
rect 4663 6780 4675 6783
rect 4890 6780 4896 6792
rect 4663 6752 4896 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4890 6740 4896 6752
rect 4948 6780 4954 6792
rect 5258 6780 5264 6792
rect 4948 6752 5264 6780
rect 4948 6740 4954 6752
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5718 6780 5724 6792
rect 5491 6752 5724 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 8168 6752 8217 6780
rect 8168 6740 8174 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8757 6783 8815 6789
rect 8757 6749 8769 6783
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 3421 6715 3479 6721
rect 3421 6712 3433 6715
rect 3384 6684 3433 6712
rect 3384 6672 3390 6684
rect 3421 6681 3433 6684
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 8496 6712 8524 6743
rect 7892 6684 8524 6712
rect 8772 6712 8800 6743
rect 8938 6712 8944 6724
rect 8772 6684 8944 6712
rect 7892 6672 7898 6684
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2188 6616 2789 6644
rect 2188 6604 2194 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3602 6644 3608 6656
rect 3099 6616 3608 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 4614 6644 4620 6656
rect 4203 6616 4620 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 7926 6644 7932 6656
rect 7791 6616 7932 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 9122 6644 9128 6656
rect 8076 6616 9128 6644
rect 8076 6604 8082 6616
rect 9122 6604 9128 6616
rect 9180 6644 9186 6656
rect 9416 6644 9444 6743
rect 9180 6616 9444 6644
rect 9180 6604 9186 6616
rect 1104 6554 9844 6576
rect 1104 6502 2702 6554
rect 2754 6502 2766 6554
rect 2818 6502 2830 6554
rect 2882 6502 2894 6554
rect 2946 6502 2958 6554
rect 3010 6502 4887 6554
rect 4939 6502 4951 6554
rect 5003 6502 5015 6554
rect 5067 6502 5079 6554
rect 5131 6502 5143 6554
rect 5195 6502 7072 6554
rect 7124 6502 7136 6554
rect 7188 6502 7200 6554
rect 7252 6502 7264 6554
rect 7316 6502 7328 6554
rect 7380 6502 9257 6554
rect 9309 6502 9321 6554
rect 9373 6502 9385 6554
rect 9437 6502 9449 6554
rect 9501 6502 9513 6554
rect 9565 6502 9844 6554
rect 1104 6480 9844 6502
rect 1946 6400 1952 6452
rect 2004 6400 2010 6452
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2406 6440 2412 6452
rect 2363 6412 2412 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6409 7251 6443
rect 7193 6403 7251 6409
rect 1854 6381 1860 6384
rect 1831 6375 1860 6381
rect 1831 6341 1843 6375
rect 1831 6335 1860 6341
rect 1854 6332 1860 6335
rect 1912 6332 1918 6384
rect 1964 6372 1992 6400
rect 2041 6375 2099 6381
rect 2041 6372 2053 6375
rect 1964 6344 2053 6372
rect 2041 6341 2053 6344
rect 2087 6341 2099 6375
rect 2041 6335 2099 6341
rect 5718 6332 5724 6384
rect 5776 6372 5782 6384
rect 5776 6344 6040 6372
rect 5776 6332 5782 6344
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 1964 6236 1992 6267
rect 2130 6264 2136 6316
rect 2188 6264 2194 6316
rect 3326 6264 3332 6316
rect 3384 6264 3390 6316
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 1820 6208 1992 6236
rect 1820 6196 1826 6208
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3200 6208 3801 6236
rect 3200 6196 3206 6208
rect 3789 6205 3801 6208
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4246 6236 4252 6248
rect 4111 6208 4252 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 5000 6236 5028 6267
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 5920 6236 5948 6267
rect 5000 6208 5948 6236
rect 6012 6236 6040 6344
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6144 6276 7021 6304
rect 6144 6264 6150 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7208 6304 7236 6403
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7208 6276 7297 6304
rect 7009 6267 7067 6273
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 7285 6267 7343 6273
rect 7576 6276 8401 6304
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 6012 6208 6377 6236
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 5000 6168 5028 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 7576 6236 7604 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8536 6276 8953 6304
rect 8536 6264 8542 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 6365 6199 6423 6205
rect 6840 6208 7604 6236
rect 1627 6140 5028 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 5258 6128 5264 6180
rect 5316 6168 5322 6180
rect 6840 6177 6868 6208
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 8168 6208 8217 6236
rect 8168 6196 8174 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 9214 6196 9220 6248
rect 9272 6196 9278 6248
rect 6825 6171 6883 6177
rect 5316 6140 6132 6168
rect 5316 6128 5322 6140
rect 3418 6060 3424 6112
rect 3476 6060 3482 6112
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5718 6100 5724 6112
rect 5123 6072 5724 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5994 6060 6000 6112
rect 6052 6060 6058 6112
rect 6104 6100 6132 6140
rect 6825 6137 6837 6171
rect 6871 6137 6883 6171
rect 6825 6131 6883 6137
rect 7466 6128 7472 6180
rect 7524 6128 7530 6180
rect 8478 6128 8484 6180
rect 8536 6128 8542 6180
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 6104 6072 7757 6100
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 1104 6010 9844 6032
rect 1104 5958 2042 6010
rect 2094 5958 2106 6010
rect 2158 5958 2170 6010
rect 2222 5958 2234 6010
rect 2286 5958 2298 6010
rect 2350 5958 4227 6010
rect 4279 5958 4291 6010
rect 4343 5958 4355 6010
rect 4407 5958 4419 6010
rect 4471 5958 4483 6010
rect 4535 5958 6412 6010
rect 6464 5958 6476 6010
rect 6528 5958 6540 6010
rect 6592 5958 6604 6010
rect 6656 5958 6668 6010
rect 6720 5958 8597 6010
rect 8649 5958 8661 6010
rect 8713 5958 8725 6010
rect 8777 5958 8789 6010
rect 8841 5958 8853 6010
rect 8905 5958 9844 6010
rect 1104 5936 9844 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 6086 5856 6092 5908
rect 6144 5856 6150 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 8938 5896 8944 5908
rect 6880 5868 8944 5896
rect 6880 5856 6886 5868
rect 8938 5856 8944 5868
rect 8996 5896 9002 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 8996 5868 9321 5896
rect 8996 5856 9002 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 4246 5788 4252 5840
rect 4304 5828 4310 5840
rect 4798 5828 4804 5840
rect 4304 5800 4804 5828
rect 4304 5788 4310 5800
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 6181 5831 6239 5837
rect 6181 5828 6193 5831
rect 5460 5800 6193 5828
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 4816 5760 4844 5788
rect 5460 5769 5488 5800
rect 6181 5797 6193 5800
rect 6227 5797 6239 5831
rect 6181 5791 6239 5797
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 8021 5831 8079 5837
rect 8021 5828 8033 5831
rect 7892 5800 8033 5828
rect 7892 5788 7898 5800
rect 8021 5797 8033 5800
rect 8067 5797 8079 5831
rect 8021 5791 8079 5797
rect 3476 5732 4568 5760
rect 3476 5720 3482 5732
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 4540 5701 4568 5732
rect 4724 5732 4844 5760
rect 5445 5763 5503 5769
rect 4724 5701 4752 5732
rect 5445 5729 5457 5763
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 5920 5732 6929 5760
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1544 5664 1869 5692
rect 1544 5652 1550 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5552 5692 5580 5720
rect 5920 5701 5948 5732
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 7650 5760 7656 5772
rect 6917 5723 6975 5729
rect 7116 5732 7656 5760
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 4847 5664 5488 5692
rect 5552 5664 5733 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 4448 5624 4476 5655
rect 4396 5596 4752 5624
rect 4396 5584 4402 5596
rect 4724 5568 4752 5596
rect 1670 5516 1676 5568
rect 1728 5516 1734 5568
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 3384 5528 4261 5556
rect 3384 5516 3390 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4249 5519 4307 5525
rect 4706 5516 4712 5568
rect 4764 5516 4770 5568
rect 5460 5556 5488 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6362 5692 6368 5704
rect 6052 5664 6368 5692
rect 6052 5652 6058 5664
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 6638 5692 6644 5704
rect 6503 5664 6644 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 6638 5652 6644 5664
rect 6696 5692 6702 5704
rect 7116 5701 7144 5732
rect 7650 5720 7656 5732
rect 7708 5760 7714 5772
rect 7708 5732 8984 5760
rect 7708 5720 7714 5732
rect 7101 5695 7159 5701
rect 6696 5664 7052 5692
rect 6696 5652 6702 5664
rect 5626 5633 5632 5636
rect 5603 5627 5632 5633
rect 5603 5593 5615 5627
rect 5603 5587 5632 5593
rect 5626 5584 5632 5587
rect 5684 5584 5690 5636
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5593 5871 5627
rect 5813 5587 5871 5593
rect 5718 5556 5724 5568
rect 5460 5528 5724 5556
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 5828 5556 5856 5587
rect 6270 5584 6276 5636
rect 6328 5624 6334 5636
rect 6733 5627 6791 5633
rect 6733 5624 6745 5627
rect 6328 5596 6745 5624
rect 6328 5584 6334 5596
rect 6733 5593 6745 5596
rect 6779 5593 6791 5627
rect 6733 5587 6791 5593
rect 6822 5584 6828 5636
rect 6880 5584 6886 5636
rect 7024 5624 7052 5664
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 7101 5655 7159 5661
rect 7208 5664 7757 5692
rect 7208 5624 7236 5664
rect 7745 5661 7757 5664
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 7883 5695 7941 5701
rect 7883 5661 7895 5695
rect 7929 5692 7941 5695
rect 8018 5692 8024 5704
rect 7929 5664 8024 5692
rect 7929 5661 7941 5664
rect 7883 5655 7941 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8956 5701 8984 5732
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8260 5664 8769 5692
rect 8260 5652 8266 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 7024 5596 7236 5624
rect 7285 5627 7343 5633
rect 7285 5593 7297 5627
rect 7331 5624 7343 5627
rect 7466 5624 7472 5636
rect 7331 5596 7472 5624
rect 7331 5593 7343 5596
rect 7285 5587 7343 5593
rect 7466 5584 7472 5596
rect 7524 5624 7530 5636
rect 9125 5627 9183 5633
rect 7524 5596 8340 5624
rect 7524 5584 7530 5596
rect 6914 5556 6920 5568
rect 5828 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 8312 5565 8340 5596
rect 9125 5593 9137 5627
rect 9171 5624 9183 5627
rect 9214 5624 9220 5636
rect 9171 5596 9220 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5525 8355 5559
rect 8297 5519 8355 5525
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9140 5556 9168 5587
rect 9214 5584 9220 5596
rect 9272 5584 9278 5636
rect 8996 5528 9168 5556
rect 8996 5516 9002 5528
rect 1104 5466 9844 5488
rect 1104 5414 2702 5466
rect 2754 5414 2766 5466
rect 2818 5414 2830 5466
rect 2882 5414 2894 5466
rect 2946 5414 2958 5466
rect 3010 5414 4887 5466
rect 4939 5414 4951 5466
rect 5003 5414 5015 5466
rect 5067 5414 5079 5466
rect 5131 5414 5143 5466
rect 5195 5414 7072 5466
rect 7124 5414 7136 5466
rect 7188 5414 7200 5466
rect 7252 5414 7264 5466
rect 7316 5414 7328 5466
rect 7380 5414 9257 5466
rect 9309 5414 9321 5466
rect 9373 5414 9385 5466
rect 9437 5414 9449 5466
rect 9501 5414 9513 5466
rect 9565 5414 9844 5466
rect 1104 5392 9844 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 1486 5352 1492 5364
rect 1443 5324 1492 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 2133 5355 2191 5361
rect 2133 5321 2145 5355
rect 2179 5321 2191 5355
rect 2133 5315 2191 5321
rect 1762 5244 1768 5296
rect 1820 5244 1826 5296
rect 1903 5287 1961 5293
rect 1903 5253 1915 5287
rect 1949 5284 1961 5287
rect 2148 5284 2176 5315
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 3108 5324 3801 5352
rect 3108 5312 3114 5324
rect 3789 5321 3801 5324
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 4856 5324 5457 5352
rect 4856 5312 4862 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5445 5315 5503 5321
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5684 5324 6377 5352
rect 5684 5312 5690 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 6972 5324 7297 5352
rect 6972 5312 6978 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 7285 5315 7343 5321
rect 1949 5256 2176 5284
rect 1949 5253 1961 5256
rect 1903 5247 1961 5253
rect 2590 5244 2596 5296
rect 2648 5284 2654 5296
rect 2685 5287 2743 5293
rect 2685 5284 2697 5287
rect 2648 5256 2697 5284
rect 2648 5244 2654 5256
rect 2685 5253 2697 5256
rect 2731 5253 2743 5287
rect 2685 5247 2743 5253
rect 2774 5244 2780 5296
rect 2832 5244 2838 5296
rect 3142 5244 3148 5296
rect 3200 5244 3206 5296
rect 3345 5287 3403 5293
rect 3345 5284 3357 5287
rect 3252 5256 3357 5284
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1688 5080 1716 5179
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 2884 5216 3096 5217
rect 3252 5216 3280 5256
rect 3345 5253 3357 5256
rect 3391 5253 3403 5287
rect 3345 5247 3403 5253
rect 5258 5244 5264 5296
rect 5316 5284 5322 5296
rect 6270 5284 6276 5296
rect 5316 5256 6276 5284
rect 5316 5244 5322 5256
rect 6270 5244 6276 5256
rect 6328 5284 6334 5296
rect 7374 5284 7380 5296
rect 6328 5256 7380 5284
rect 6328 5244 6334 5256
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 2464 5189 3280 5216
rect 2464 5188 2912 5189
rect 3068 5188 3280 5189
rect 4249 5219 4307 5225
rect 2464 5176 2470 5188
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4338 5216 4344 5228
rect 4295 5188 4344 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4706 5216 4712 5228
rect 4479 5188 4712 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4856 5188 4997 5216
rect 4856 5176 4862 5188
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5592 5188 5733 5216
rect 5592 5176 5598 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6236 5188 6561 5216
rect 6236 5176 6242 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6730 5176 6736 5228
rect 6788 5176 6794 5228
rect 7190 5176 7196 5228
rect 7248 5176 7254 5228
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 2041 5151 2099 5157
rect 2041 5148 2053 5151
rect 1912 5120 2053 5148
rect 1912 5108 1918 5120
rect 2041 5117 2053 5120
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2498 5148 2504 5160
rect 2363 5120 2504 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2498 5108 2504 5120
rect 2556 5148 2562 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 2556 5120 4905 5148
rect 2556 5108 2562 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 1946 5080 1952 5092
rect 1688 5052 1952 5080
rect 1946 5040 1952 5052
rect 2004 5040 2010 5092
rect 4522 5040 4528 5092
rect 4580 5080 4586 5092
rect 4617 5083 4675 5089
rect 4617 5080 4629 5083
rect 4580 5052 4629 5080
rect 4580 5040 4586 5052
rect 4617 5049 4629 5052
rect 4663 5049 4675 5083
rect 4908 5080 4936 5111
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 5626 5108 5632 5160
rect 5684 5108 5690 5160
rect 5810 5108 5816 5160
rect 5868 5108 5874 5160
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 7009 5083 7067 5089
rect 4908 5052 6408 5080
rect 4617 5043 4675 5049
rect 6380 5024 6408 5052
rect 7009 5049 7021 5083
rect 7055 5080 7067 5083
rect 7300 5080 7328 5179
rect 7466 5176 7472 5228
rect 7524 5176 7530 5228
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8386 5216 8392 5228
rect 8076 5188 8392 5216
rect 8076 5176 8082 5188
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 7650 5080 7656 5092
rect 7055 5052 7656 5080
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 8202 5040 8208 5092
rect 8260 5040 8266 5092
rect 3326 4972 3332 5024
rect 3384 4972 3390 5024
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 3694 5012 3700 5024
rect 3559 4984 3700 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4246 5012 4252 5024
rect 4111 4984 4252 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4709 5015 4767 5021
rect 4709 4981 4721 5015
rect 4755 5012 4767 5015
rect 4982 5012 4988 5024
rect 4755 4984 4988 5012
rect 4755 4981 4767 4984
rect 4709 4975 4767 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 7742 5012 7748 5024
rect 6420 4984 7748 5012
rect 6420 4972 6426 4984
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 1104 4922 9844 4944
rect 1104 4870 2042 4922
rect 2094 4870 2106 4922
rect 2158 4870 2170 4922
rect 2222 4870 2234 4922
rect 2286 4870 2298 4922
rect 2350 4870 4227 4922
rect 4279 4870 4291 4922
rect 4343 4870 4355 4922
rect 4407 4870 4419 4922
rect 4471 4870 4483 4922
rect 4535 4870 6412 4922
rect 6464 4870 6476 4922
rect 6528 4870 6540 4922
rect 6592 4870 6604 4922
rect 6656 4870 6668 4922
rect 6720 4870 8597 4922
rect 8649 4870 8661 4922
rect 8713 4870 8725 4922
rect 8777 4870 8789 4922
rect 8841 4870 8853 4922
rect 8905 4870 9844 4922
rect 1104 4848 9844 4870
rect 1210 4768 1216 4820
rect 1268 4808 1274 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1268 4780 1501 4808
rect 1268 4768 1274 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1489 4771 1547 4777
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 1854 4808 1860 4820
rect 1811 4780 1860 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2832 4780 2881 4808
rect 2832 4768 2838 4780
rect 2869 4777 2881 4780
rect 2915 4808 2927 4811
rect 3786 4808 3792 4820
rect 2915 4780 3792 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 5902 4808 5908 4820
rect 5215 4780 5908 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8352 4780 8524 4808
rect 8352 4768 8358 4780
rect 6178 4740 6184 4752
rect 1964 4712 6184 4740
rect 1670 4564 1676 4616
rect 1728 4564 1734 4616
rect 1302 4496 1308 4548
rect 1360 4536 1366 4548
rect 1964 4545 1992 4712
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 4249 4675 4307 4681
rect 3752 4644 4016 4672
rect 3752 4632 3758 4644
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3200 4576 3249 4604
rect 3200 4564 3206 4576
rect 3237 4573 3249 4576
rect 3283 4604 3295 4607
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 3283 4576 3341 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 1949 4539 2007 4545
rect 1949 4536 1961 4539
rect 1360 4508 1961 4536
rect 1360 4496 1366 4508
rect 1949 4505 1961 4508
rect 1995 4505 2007 4539
rect 1949 4499 2007 4505
rect 2133 4539 2191 4545
rect 2133 4505 2145 4539
rect 2179 4536 2191 4539
rect 2406 4536 2412 4548
rect 2179 4508 2412 4536
rect 2179 4505 2191 4508
rect 2133 4499 2191 4505
rect 2406 4496 2412 4508
rect 2464 4536 2470 4548
rect 2464 4508 2774 4536
rect 2464 4496 2470 4508
rect 2746 4468 2774 4508
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 3528 4536 3556 4567
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3988 4604 4016 4644
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4614 4672 4620 4684
rect 4295 4644 4620 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4724 4681 4752 4712
rect 6178 4700 6184 4712
rect 6236 4700 6242 4752
rect 6733 4743 6791 4749
rect 6733 4709 6745 4743
rect 6779 4740 6791 4743
rect 6914 4740 6920 4752
rect 6779 4712 6920 4740
rect 6779 4709 6791 4712
rect 6733 4703 6791 4709
rect 6914 4700 6920 4712
rect 6972 4740 6978 4752
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 6972 4712 7481 4740
rect 6972 4700 6978 4712
rect 7469 4709 7481 4712
rect 7515 4740 7527 4743
rect 8018 4740 8024 4752
rect 7515 4712 8024 4740
rect 7515 4709 7527 4712
rect 7469 4703 7527 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 8496 4749 8524 4780
rect 8481 4743 8539 4749
rect 8481 4709 8493 4743
rect 8527 4709 8539 4743
rect 8481 4703 8539 4709
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4641 4767 4675
rect 8294 4672 8300 4684
rect 4709 4635 4767 4641
rect 6564 4644 8300 4672
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 3988 4576 4353 4604
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 6564 4613 6592 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6972 4576 7021 4604
rect 6972 4564 6978 4576
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7285 4607 7343 4613
rect 7055 4576 7236 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 3108 4508 3556 4536
rect 3108 4496 3114 4508
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 7101 4539 7159 4545
rect 7101 4536 7113 4539
rect 6696 4508 7113 4536
rect 6696 4496 6702 4508
rect 7101 4505 7113 4508
rect 7147 4505 7159 4539
rect 7208 4536 7236 4576
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7374 4604 7380 4616
rect 7331 4576 7380 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7576 4536 7604 4567
rect 7650 4564 7656 4616
rect 7708 4564 7714 4616
rect 8202 4564 8208 4616
rect 8260 4564 8266 4616
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 9122 4564 9128 4616
rect 9180 4564 9186 4616
rect 7208 4508 7604 4536
rect 7101 4499 7159 4505
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 7800 4508 8953 4536
rect 7800 4496 7806 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2746 4440 3433 4468
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4614 4468 4620 4480
rect 4019 4440 4620 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 6917 4471 6975 4477
rect 6917 4468 6929 4471
rect 6880 4440 6929 4468
rect 6880 4428 6886 4440
rect 6917 4437 6929 4440
rect 6963 4437 6975 4471
rect 6917 4431 6975 4437
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9140 4468 9168 4564
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 9674 4536 9680 4548
rect 9539 4508 9680 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 8260 4440 9168 4468
rect 8260 4428 8266 4440
rect 1104 4378 9844 4400
rect 1104 4326 2702 4378
rect 2754 4326 2766 4378
rect 2818 4326 2830 4378
rect 2882 4326 2894 4378
rect 2946 4326 2958 4378
rect 3010 4326 4887 4378
rect 4939 4326 4951 4378
rect 5003 4326 5015 4378
rect 5067 4326 5079 4378
rect 5131 4326 5143 4378
rect 5195 4326 7072 4378
rect 7124 4326 7136 4378
rect 7188 4326 7200 4378
rect 7252 4326 7264 4378
rect 7316 4326 7328 4378
rect 7380 4326 9257 4378
rect 9309 4326 9321 4378
rect 9373 4326 9385 4378
rect 9437 4326 9449 4378
rect 9501 4326 9513 4378
rect 9565 4326 9844 4378
rect 1104 4304 9844 4326
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6733 4267 6791 4273
rect 6733 4264 6745 4267
rect 6236 4236 6745 4264
rect 6236 4224 6242 4236
rect 6733 4233 6745 4236
rect 6779 4233 6791 4267
rect 6733 4227 6791 4233
rect 5442 4196 5448 4208
rect 4908 4168 5448 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4908 4128 4936 4168
rect 5442 4156 5448 4168
rect 5500 4156 5506 4208
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 7650 4196 7656 4208
rect 6880 4168 6960 4196
rect 6880 4156 6886 4168
rect 4663 4100 4936 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4982 4088 4988 4140
rect 5040 4088 5046 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5258 4128 5264 4140
rect 5215 4100 5264 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 5184 4060 5212 4091
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 4939 4032 5212 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 6638 4020 6644 4072
rect 6696 4060 6702 4072
rect 6932 4069 6960 4168
rect 7392 4168 7656 4196
rect 7392 4137 7420 4168
rect 7650 4156 7656 4168
rect 7708 4156 7714 4208
rect 8110 4156 8116 4208
rect 8168 4156 8174 4208
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 8128 4128 8156 4156
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8128 4100 8585 4128
rect 7561 4091 7619 4097
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9582 4128 9588 4140
rect 9447 4100 9588 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6696 4032 6837 4060
rect 6696 4020 6702 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 4801 3995 4859 4001
rect 4801 3961 4813 3995
rect 4847 3992 4859 3995
rect 5626 3992 5632 4004
rect 4847 3964 5632 3992
rect 4847 3961 4859 3964
rect 4801 3955 4859 3961
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7469 3995 7527 4001
rect 7469 3992 7481 3995
rect 6788 3964 7481 3992
rect 6788 3952 6794 3964
rect 7469 3961 7481 3964
rect 7515 3961 7527 3995
rect 7576 3992 7604 4091
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7708 4032 7849 4060
rect 7708 4020 7714 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 7926 4020 7932 4072
rect 7984 4020 7990 4072
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4060 8171 4063
rect 8202 4060 8208 4072
rect 8159 4032 8208 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 9674 4060 9680 4072
rect 8352 4032 9680 4060
rect 8352 4020 8358 4032
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 7576 3964 8248 3992
rect 7469 3955 7527 3961
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2866 3924 2872 3936
rect 1627 3896 2872 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2866 3884 2872 3896
rect 2924 3924 2930 3936
rect 3142 3924 3148 3936
rect 2924 3896 3148 3924
rect 2924 3884 2930 3896
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4120 3896 4721 3924
rect 4120 3884 4126 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4948 3896 5089 3924
rect 4948 3884 4954 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6328 3896 6377 3924
rect 6328 3884 6334 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 7653 3927 7711 3933
rect 7653 3924 7665 3927
rect 7616 3896 7665 3924
rect 7616 3884 7622 3896
rect 7653 3893 7665 3896
rect 7699 3893 7711 3927
rect 8220 3924 8248 3964
rect 8938 3924 8944 3936
rect 8220 3896 8944 3924
rect 7653 3887 7711 3893
rect 8938 3884 8944 3896
rect 8996 3924 9002 3936
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 8996 3896 9229 3924
rect 8996 3884 9002 3896
rect 9217 3893 9229 3896
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 1104 3834 9844 3856
rect 1104 3782 2042 3834
rect 2094 3782 2106 3834
rect 2158 3782 2170 3834
rect 2222 3782 2234 3834
rect 2286 3782 2298 3834
rect 2350 3782 4227 3834
rect 4279 3782 4291 3834
rect 4343 3782 4355 3834
rect 4407 3782 4419 3834
rect 4471 3782 4483 3834
rect 4535 3782 6412 3834
rect 6464 3782 6476 3834
rect 6528 3782 6540 3834
rect 6592 3782 6604 3834
rect 6656 3782 6668 3834
rect 6720 3782 8597 3834
rect 8649 3782 8661 3834
rect 8713 3782 8725 3834
rect 8777 3782 8789 3834
rect 8841 3782 8853 3834
rect 8905 3782 9844 3834
rect 1104 3760 9844 3782
rect 1578 3680 1584 3732
rect 1636 3720 1642 3732
rect 1857 3723 1915 3729
rect 1857 3720 1869 3723
rect 1636 3692 1869 3720
rect 1636 3680 1642 3692
rect 1857 3689 1869 3692
rect 1903 3689 1915 3723
rect 1857 3683 1915 3689
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 2096 3692 2513 3720
rect 2096 3680 2102 3692
rect 2501 3689 2513 3692
rect 2547 3720 2559 3723
rect 2777 3723 2835 3729
rect 2547 3692 2636 3720
rect 2547 3689 2559 3692
rect 2501 3683 2559 3689
rect 2608 3661 2636 3692
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3326 3720 3332 3732
rect 2823 3692 3332 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 4246 3720 4252 3732
rect 3651 3692 4252 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 4246 3680 4252 3692
rect 4304 3720 4310 3732
rect 4709 3723 4767 3729
rect 4709 3720 4721 3723
rect 4304 3692 4721 3720
rect 4304 3680 4310 3692
rect 4709 3689 4721 3692
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 5350 3680 5356 3732
rect 5408 3680 5414 3732
rect 5905 3723 5963 3729
rect 5905 3689 5917 3723
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 1949 3655 2007 3661
rect 1949 3621 1961 3655
rect 1995 3652 2007 3655
rect 2593 3655 2651 3661
rect 1995 3624 2544 3652
rect 1995 3621 2007 3624
rect 1949 3615 2007 3621
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 1811 3556 2421 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2409 3553 2421 3556
rect 2455 3553 2467 3587
rect 2409 3547 2467 3553
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 2424 3448 2452 3547
rect 2516 3528 2544 3624
rect 2593 3621 2605 3655
rect 2639 3621 2651 3655
rect 2593 3615 2651 3621
rect 2608 3584 2636 3615
rect 3234 3612 3240 3664
rect 3292 3612 3298 3664
rect 4893 3655 4951 3661
rect 4893 3621 4905 3655
rect 4939 3652 4951 3655
rect 5920 3652 5948 3683
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 6328 3692 6653 3720
rect 6328 3680 6334 3692
rect 6641 3689 6653 3692
rect 6687 3689 6699 3723
rect 6641 3683 6699 3689
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 4939 3624 5856 3652
rect 5920 3624 9045 3652
rect 4939 3621 4951 3624
rect 4893 3615 4951 3621
rect 3252 3584 3280 3612
rect 3510 3584 3516 3596
rect 2608 3556 3188 3584
rect 3252 3556 3516 3584
rect 2498 3476 2504 3528
rect 2556 3476 2562 3528
rect 3160 3525 3188 3556
rect 3510 3544 3516 3556
rect 3568 3584 3574 3596
rect 5718 3584 5724 3596
rect 3568 3556 4292 3584
rect 3568 3544 3574 3556
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 2866 3448 2872 3460
rect 2424 3420 2872 3448
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 2961 3451 3019 3457
rect 2961 3417 2973 3451
rect 3007 3417 3019 3451
rect 3068 3448 3096 3479
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3292 3488 3341 3516
rect 3292 3476 3298 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3467 3488 3801 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4264 3525 4292 3556
rect 4448 3556 5724 3584
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4448 3448 4476 3556
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5828 3593 5856 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9033 3615 9091 3621
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3553 5871 3587
rect 7558 3584 7564 3596
rect 5813 3547 5871 3553
rect 6932 3556 7564 3584
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5258 3516 5264 3528
rect 5031 3488 5264 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5408 3488 5549 3516
rect 5408 3476 5414 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5736 3516 5764 3544
rect 6178 3516 6184 3528
rect 5736 3488 6184 3516
rect 5537 3479 5595 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6932 3525 6960 3556
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 8444 3556 8493 3584
rect 8444 3544 8450 3556
rect 8481 3553 8493 3556
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 9674 3584 9680 3596
rect 9539 3556 9680 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7147 3488 7297 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 3068 3420 4476 3448
rect 4525 3451 4583 3457
rect 2961 3411 3019 3417
rect 4525 3417 4537 3451
rect 4571 3448 4583 3451
rect 4614 3448 4620 3460
rect 4571 3420 4620 3448
rect 4571 3417 4583 3420
rect 4525 3411 4583 3417
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 2004 3352 2145 3380
rect 2004 3340 2010 3352
rect 2133 3349 2145 3352
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 2751 3383 2809 3389
rect 2751 3380 2763 3383
rect 2648 3352 2763 3380
rect 2648 3340 2654 3352
rect 2751 3349 2763 3352
rect 2797 3349 2809 3383
rect 2976 3380 3004 3411
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 4741 3451 4799 3457
rect 4741 3417 4753 3451
rect 4787 3448 4799 3451
rect 4890 3448 4896 3460
rect 4787 3420 4896 3448
rect 4787 3417 4799 3420
rect 4741 3411 4799 3417
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 5169 3451 5227 3457
rect 5169 3417 5181 3451
rect 5215 3417 5227 3451
rect 6196 3448 6224 3476
rect 7190 3448 7196 3460
rect 6196 3420 7196 3448
rect 5169 3411 5227 3417
rect 3050 3380 3056 3392
rect 2976 3352 3056 3380
rect 2751 3343 2809 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 4157 3383 4215 3389
rect 4157 3380 4169 3383
rect 3384 3352 4169 3380
rect 3384 3340 3390 3352
rect 4157 3349 4169 3352
rect 4203 3349 4215 3383
rect 4157 3343 4215 3349
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 4982 3380 4988 3392
rect 4488 3352 4988 3380
rect 4488 3340 4494 3352
rect 4982 3340 4988 3352
rect 5040 3380 5046 3392
rect 5184 3380 5212 3411
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 7300 3448 7328 3479
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 7834 3516 7840 3528
rect 7699 3488 7840 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8182 3519 8240 3525
rect 8182 3485 8194 3519
rect 8228 3516 8240 3519
rect 8294 3516 8300 3528
rect 8228 3488 8300 3516
rect 8228 3485 8240 3488
rect 8182 3479 8240 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 7466 3448 7472 3460
rect 7300 3420 7472 3448
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 9030 3448 9036 3460
rect 7616 3420 9036 3448
rect 7616 3408 7622 3420
rect 8128 3392 8156 3420
rect 9030 3408 9036 3420
rect 9088 3408 9094 3460
rect 5040 3352 5212 3380
rect 5040 3340 5046 3352
rect 6086 3340 6092 3392
rect 6144 3340 6150 3392
rect 6825 3383 6883 3389
rect 6825 3349 6837 3383
rect 6871 3380 6883 3383
rect 7742 3380 7748 3392
rect 6871 3352 7748 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8110 3340 8116 3392
rect 8168 3340 8174 3392
rect 1104 3290 9844 3312
rect 1104 3238 2702 3290
rect 2754 3238 2766 3290
rect 2818 3238 2830 3290
rect 2882 3238 2894 3290
rect 2946 3238 2958 3290
rect 3010 3238 4887 3290
rect 4939 3238 4951 3290
rect 5003 3238 5015 3290
rect 5067 3238 5079 3290
rect 5131 3238 5143 3290
rect 5195 3238 7072 3290
rect 7124 3238 7136 3290
rect 7188 3238 7200 3290
rect 7252 3238 7264 3290
rect 7316 3238 7328 3290
rect 7380 3238 9257 3290
rect 9309 3238 9321 3290
rect 9373 3238 9385 3290
rect 9437 3238 9449 3290
rect 9501 3238 9513 3290
rect 9565 3238 9844 3290
rect 1104 3216 9844 3238
rect 3234 3136 3240 3188
rect 3292 3136 3298 3188
rect 4246 3136 4252 3188
rect 4304 3136 4310 3188
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 5442 3176 5448 3188
rect 4939 3148 5448 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 2869 3111 2927 3117
rect 2869 3077 2881 3111
rect 2915 3108 2927 3111
rect 3326 3108 3332 3120
rect 2915 3080 3332 3108
rect 2915 3077 2927 3080
rect 2869 3071 2927 3077
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 4525 3111 4583 3117
rect 4525 3108 4537 3111
rect 4172 3080 4537 3108
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 2774 3040 2780 3052
rect 2731 3012 2780 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 2961 3003 3019 3009
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2976 2972 3004 3003
rect 3142 3000 3148 3052
rect 3200 3000 3206 3052
rect 4172 3049 4200 3080
rect 4525 3077 4537 3080
rect 4571 3108 4583 3111
rect 4614 3108 4620 3120
rect 4571 3080 4620 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 4755 3077 4813 3083
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4755 3043 4767 3077
rect 4801 3074 4813 3077
rect 4801 3052 4855 3074
rect 4801 3043 4804 3052
rect 4755 3040 4804 3043
rect 4488 3012 4804 3040
rect 4488 3000 4494 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 5000 3049 5028 3148
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6144 3148 7021 3176
rect 6144 3136 6150 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7009 3139 7067 3145
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7561 3179 7619 3185
rect 7561 3176 7573 3179
rect 7524 3148 7573 3176
rect 7524 3136 7530 3148
rect 7561 3145 7573 3148
rect 7607 3145 7619 3179
rect 7561 3139 7619 3145
rect 7834 3136 7840 3188
rect 7892 3136 7898 3188
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 7984 3148 9137 3176
rect 7984 3136 7990 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9125 3139 9183 3145
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5258 3000 5264 3052
rect 5316 3000 5322 3052
rect 5460 3040 5488 3136
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 5810 3108 5816 3120
rect 5767 3080 5816 3108
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 5810 3068 5816 3080
rect 5868 3108 5874 3120
rect 8757 3111 8815 3117
rect 8757 3108 8769 3111
rect 5868 3080 6684 3108
rect 5868 3068 5874 3080
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5460 3012 6009 3040
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6178 3000 6184 3052
rect 6236 3000 6242 3052
rect 6656 3049 6684 3080
rect 7760 3080 8769 3108
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7466 3040 7472 3052
rect 7239 3012 7472 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 3510 2972 3516 2984
rect 2648 2944 3516 2972
rect 2648 2932 2654 2944
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 4172 2944 5089 2972
rect 4172 2916 4200 2944
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 6089 2975 6147 2981
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6135 2944 6561 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 7576 2972 7604 3003
rect 7650 3000 7656 3052
rect 7708 3040 7714 3052
rect 7760 3049 7788 3080
rect 8757 3077 8769 3080
rect 8803 3077 8815 3111
rect 8757 3071 8815 3077
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7708 3012 7757 3040
rect 7708 3000 7714 3012
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8018 2972 8024 2984
rect 7576 2944 8024 2972
rect 6549 2935 6607 2941
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8404 2972 8432 3003
rect 8570 3000 8576 3052
rect 8628 3000 8634 3052
rect 8772 3040 8800 3071
rect 9030 3068 9036 3120
rect 9088 3068 9094 3120
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8772 3012 8953 3040
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 8352 2944 8432 2972
rect 8496 2944 9413 2972
rect 8352 2932 8358 2944
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 2556 2876 2697 2904
rect 2556 2864 2562 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 2685 2867 2743 2873
rect 4154 2864 4160 2916
rect 4212 2864 4218 2916
rect 4246 2864 4252 2916
rect 4304 2904 4310 2916
rect 4304 2876 4752 2904
rect 4304 2864 4310 2876
rect 4172 2836 4200 2864
rect 4724 2845 4752 2876
rect 6914 2864 6920 2916
rect 6972 2904 6978 2916
rect 7834 2904 7840 2916
rect 6972 2876 7840 2904
rect 6972 2864 6978 2876
rect 7834 2864 7840 2876
rect 7892 2904 7898 2916
rect 7929 2907 7987 2913
rect 7929 2904 7941 2907
rect 7892 2876 7941 2904
rect 7892 2864 7898 2876
rect 7929 2873 7941 2876
rect 7975 2873 7987 2907
rect 8036 2904 8064 2932
rect 8496 2904 8524 2944
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9401 2935 9459 2941
rect 8036 2876 8524 2904
rect 7929 2867 7987 2873
rect 4433 2839 4491 2845
rect 4433 2836 4445 2839
rect 4172 2808 4445 2836
rect 4433 2805 4445 2808
rect 4479 2805 4491 2839
rect 4433 2799 4491 2805
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2805 4767 2839
rect 4709 2799 4767 2805
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6328 2808 6377 2836
rect 6328 2796 6334 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 7944 2836 7972 2867
rect 8570 2836 8576 2848
rect 7944 2808 8576 2836
rect 6365 2799 6423 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 1104 2746 9844 2768
rect 1104 2694 2042 2746
rect 2094 2694 2106 2746
rect 2158 2694 2170 2746
rect 2222 2694 2234 2746
rect 2286 2694 2298 2746
rect 2350 2694 4227 2746
rect 4279 2694 4291 2746
rect 4343 2694 4355 2746
rect 4407 2694 4419 2746
rect 4471 2694 4483 2746
rect 4535 2694 6412 2746
rect 6464 2694 6476 2746
rect 6528 2694 6540 2746
rect 6592 2694 6604 2746
rect 6656 2694 6668 2746
rect 6720 2694 8597 2746
rect 8649 2694 8661 2746
rect 8713 2694 8725 2746
rect 8777 2694 8789 2746
rect 8841 2694 8853 2746
rect 8905 2694 9844 2746
rect 1104 2672 9844 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3050 2632 3056 2644
rect 2832 2604 3056 2632
rect 2832 2592 2838 2604
rect 3050 2592 3056 2604
rect 3108 2632 3114 2644
rect 3513 2635 3571 2641
rect 3513 2632 3525 2635
rect 3108 2604 3525 2632
rect 3108 2592 3114 2604
rect 3513 2601 3525 2604
rect 3559 2632 3571 2635
rect 3970 2632 3976 2644
rect 3559 2604 3976 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4798 2632 4804 2644
rect 4203 2604 4804 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5258 2592 5264 2644
rect 5316 2632 5322 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 5316 2604 5457 2632
rect 5316 2592 5322 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 5445 2595 5503 2601
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8018 2632 8024 2644
rect 7975 2604 8024 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8294 2592 8300 2644
rect 8352 2592 8358 2644
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8536 2604 8677 2632
rect 8536 2592 8542 2604
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 8665 2595 8723 2601
rect 8312 2496 8340 2592
rect 8036 2468 8340 2496
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 5316 2400 5641 2428
rect 5316 2388 5322 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 6328 2400 6469 2428
rect 6328 2388 6334 2400
rect 6457 2397 6469 2400
rect 6503 2397 6515 2431
rect 6457 2391 6515 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7515 2400 7604 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 5077 2363 5135 2369
rect 5077 2360 5089 2363
rect 4580 2332 5089 2360
rect 4580 2320 4586 2332
rect 5077 2329 5089 2332
rect 5123 2329 5135 2363
rect 5077 2323 5135 2329
rect 5810 2320 5816 2372
rect 5868 2360 5874 2372
rect 6825 2363 6883 2369
rect 6825 2360 6837 2363
rect 5868 2332 6837 2360
rect 5868 2320 5874 2332
rect 6825 2329 6837 2332
rect 6871 2329 6883 2363
rect 6825 2323 6883 2329
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7576 2301 7604 2400
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8036 2437 8064 2468
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8128 2360 8156 2391
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8444 2400 8493 2428
rect 8444 2388 8450 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 7760 2332 8156 2360
rect 7760 2304 7788 2332
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 6972 2264 7297 2292
rect 6972 2252 6978 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 7561 2295 7619 2301
rect 7561 2261 7573 2295
rect 7607 2261 7619 2295
rect 7561 2255 7619 2261
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 1104 2202 9844 2224
rect 1104 2150 2702 2202
rect 2754 2150 2766 2202
rect 2818 2150 2830 2202
rect 2882 2150 2894 2202
rect 2946 2150 2958 2202
rect 3010 2150 4887 2202
rect 4939 2150 4951 2202
rect 5003 2150 5015 2202
rect 5067 2150 5079 2202
rect 5131 2150 5143 2202
rect 5195 2150 7072 2202
rect 7124 2150 7136 2202
rect 7188 2150 7200 2202
rect 7252 2150 7264 2202
rect 7316 2150 7328 2202
rect 7380 2150 9257 2202
rect 9309 2150 9321 2202
rect 9373 2150 9385 2202
rect 9437 2150 9449 2202
rect 9501 2150 9513 2202
rect 9565 2150 9844 2202
rect 1104 2128 9844 2150
<< via1 >>
rect 2702 10854 2754 10906
rect 2766 10854 2818 10906
rect 2830 10854 2882 10906
rect 2894 10854 2946 10906
rect 2958 10854 3010 10906
rect 4887 10854 4939 10906
rect 4951 10854 5003 10906
rect 5015 10854 5067 10906
rect 5079 10854 5131 10906
rect 5143 10854 5195 10906
rect 7072 10854 7124 10906
rect 7136 10854 7188 10906
rect 7200 10854 7252 10906
rect 7264 10854 7316 10906
rect 7328 10854 7380 10906
rect 9257 10854 9309 10906
rect 9321 10854 9373 10906
rect 9385 10854 9437 10906
rect 9449 10854 9501 10906
rect 9513 10854 9565 10906
rect 3424 10795 3476 10804
rect 3424 10761 3441 10795
rect 3441 10761 3476 10795
rect 3424 10752 3476 10761
rect 5264 10752 5316 10804
rect 3700 10684 3752 10736
rect 3976 10684 4028 10736
rect 3608 10548 3660 10600
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 7748 10684 7800 10736
rect 5816 10616 5868 10668
rect 6092 10616 6144 10668
rect 6552 10616 6604 10668
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 4620 10548 4672 10600
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 7932 10548 7984 10600
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 6920 10480 6972 10532
rect 8116 10480 8168 10532
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3976 10412 4028 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 7012 10412 7064 10464
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 2042 10310 2094 10362
rect 2106 10310 2158 10362
rect 2170 10310 2222 10362
rect 2234 10310 2286 10362
rect 2298 10310 2350 10362
rect 4227 10310 4279 10362
rect 4291 10310 4343 10362
rect 4355 10310 4407 10362
rect 4419 10310 4471 10362
rect 4483 10310 4535 10362
rect 6412 10310 6464 10362
rect 6476 10310 6528 10362
rect 6540 10310 6592 10362
rect 6604 10310 6656 10362
rect 6668 10310 6720 10362
rect 8597 10310 8649 10362
rect 8661 10310 8713 10362
rect 8725 10310 8777 10362
rect 8789 10310 8841 10362
rect 8853 10310 8905 10362
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 5264 10140 5316 10192
rect 3608 10115 3660 10124
rect 3608 10081 3617 10115
rect 3617 10081 3651 10115
rect 3651 10081 3660 10115
rect 3608 10072 3660 10081
rect 3700 10072 3752 10124
rect 4528 10072 4580 10124
rect 5356 10072 5408 10124
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 7932 10072 7984 10124
rect 8392 10072 8444 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3976 10004 4028 10056
rect 4160 10004 4212 10056
rect 4804 10004 4856 10056
rect 6000 10004 6052 10056
rect 7012 10004 7064 10056
rect 7472 10004 7524 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 6736 9936 6788 9988
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 8392 9936 8444 9988
rect 9128 9936 9180 9988
rect 2596 9868 2648 9920
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 6276 9868 6328 9877
rect 8668 9868 8720 9920
rect 2702 9766 2754 9818
rect 2766 9766 2818 9818
rect 2830 9766 2882 9818
rect 2894 9766 2946 9818
rect 2958 9766 3010 9818
rect 4887 9766 4939 9818
rect 4951 9766 5003 9818
rect 5015 9766 5067 9818
rect 5079 9766 5131 9818
rect 5143 9766 5195 9818
rect 7072 9766 7124 9818
rect 7136 9766 7188 9818
rect 7200 9766 7252 9818
rect 7264 9766 7316 9818
rect 7328 9766 7380 9818
rect 9257 9766 9309 9818
rect 9321 9766 9373 9818
rect 9385 9766 9437 9818
rect 9449 9766 9501 9818
rect 9513 9766 9565 9818
rect 3424 9664 3476 9716
rect 7748 9664 7800 9716
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 8484 9664 8536 9716
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4068 9528 4120 9580
rect 4528 9528 4580 9580
rect 4804 9596 4856 9648
rect 6276 9596 6328 9648
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 6736 9528 6788 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 8116 9639 8168 9648
rect 8116 9605 8151 9639
rect 8151 9605 8168 9639
rect 8116 9596 8168 9605
rect 7472 9528 7524 9580
rect 7748 9528 7800 9580
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 5080 9392 5132 9444
rect 6184 9392 6236 9444
rect 7656 9460 7708 9512
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 9128 9596 9180 9648
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 6828 9435 6880 9444
rect 6828 9401 6837 9435
rect 6837 9401 6871 9435
rect 6871 9401 6880 9435
rect 6828 9392 6880 9401
rect 7472 9392 7524 9444
rect 8024 9392 8076 9444
rect 8208 9392 8260 9444
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 5448 9324 5500 9376
rect 7748 9324 7800 9376
rect 8116 9324 8168 9376
rect 9588 9324 9640 9376
rect 2042 9222 2094 9274
rect 2106 9222 2158 9274
rect 2170 9222 2222 9274
rect 2234 9222 2286 9274
rect 2298 9222 2350 9274
rect 4227 9222 4279 9274
rect 4291 9222 4343 9274
rect 4355 9222 4407 9274
rect 4419 9222 4471 9274
rect 4483 9222 4535 9274
rect 6412 9222 6464 9274
rect 6476 9222 6528 9274
rect 6540 9222 6592 9274
rect 6604 9222 6656 9274
rect 6668 9222 6720 9274
rect 8597 9222 8649 9274
rect 8661 9222 8713 9274
rect 8725 9222 8777 9274
rect 8789 9222 8841 9274
rect 8853 9222 8905 9274
rect 4620 9120 4672 9172
rect 848 9052 900 9104
rect 2412 9052 2464 9104
rect 2504 9052 2556 9104
rect 4896 9052 4948 9104
rect 7564 9052 7616 9104
rect 1860 8984 1912 9036
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 2596 8984 2648 9036
rect 5816 8984 5868 9036
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 1952 8891 2004 8900
rect 1952 8857 1969 8891
rect 1969 8857 2004 8891
rect 1952 8848 2004 8857
rect 2964 8848 3016 8900
rect 3332 8848 3384 8900
rect 4804 8916 4856 8968
rect 5724 8916 5776 8968
rect 7840 8916 7892 8968
rect 8576 8984 8628 9036
rect 9312 8984 9364 9036
rect 8392 8959 8444 8968
rect 8392 8925 8401 8959
rect 8401 8925 8435 8959
rect 8435 8925 8444 8959
rect 8392 8916 8444 8925
rect 8484 8959 8536 8968
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9036 8916 9088 8968
rect 9220 8916 9272 8968
rect 3792 8780 3844 8832
rect 5080 8780 5132 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 8208 8780 8260 8832
rect 2702 8678 2754 8730
rect 2766 8678 2818 8730
rect 2830 8678 2882 8730
rect 2894 8678 2946 8730
rect 2958 8678 3010 8730
rect 4887 8678 4939 8730
rect 4951 8678 5003 8730
rect 5015 8678 5067 8730
rect 5079 8678 5131 8730
rect 5143 8678 5195 8730
rect 7072 8678 7124 8730
rect 7136 8678 7188 8730
rect 7200 8678 7252 8730
rect 7264 8678 7316 8730
rect 7328 8678 7380 8730
rect 9257 8678 9309 8730
rect 9321 8678 9373 8730
rect 9385 8678 9437 8730
rect 9449 8678 9501 8730
rect 9513 8678 9565 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 1952 8576 2004 8628
rect 7472 8576 7524 8628
rect 8116 8576 8168 8628
rect 1308 8440 1360 8492
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 2596 8372 2648 8424
rect 4804 8508 4856 8560
rect 4712 8440 4764 8492
rect 6828 8508 6880 8560
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 4804 8372 4856 8424
rect 5080 8372 5132 8424
rect 5540 8372 5592 8424
rect 5816 8440 5868 8492
rect 6276 8440 6328 8492
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6184 8372 6236 8424
rect 6000 8304 6052 8356
rect 7012 8440 7064 8492
rect 7380 8440 7432 8492
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8576 8576 8628 8628
rect 8300 8508 8352 8560
rect 8392 8508 8444 8560
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 7104 8304 7156 8356
rect 5172 8236 5224 8288
rect 5448 8236 5500 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 5632 8236 5684 8288
rect 6552 8236 6604 8288
rect 8300 8304 8352 8356
rect 8484 8347 8536 8356
rect 8484 8313 8493 8347
rect 8493 8313 8527 8347
rect 8527 8313 8536 8347
rect 8484 8304 8536 8313
rect 9036 8236 9088 8288
rect 2042 8134 2094 8186
rect 2106 8134 2158 8186
rect 2170 8134 2222 8186
rect 2234 8134 2286 8186
rect 2298 8134 2350 8186
rect 4227 8134 4279 8186
rect 4291 8134 4343 8186
rect 4355 8134 4407 8186
rect 4419 8134 4471 8186
rect 4483 8134 4535 8186
rect 6412 8134 6464 8186
rect 6476 8134 6528 8186
rect 6540 8134 6592 8186
rect 6604 8134 6656 8186
rect 6668 8134 6720 8186
rect 8597 8134 8649 8186
rect 8661 8134 8713 8186
rect 8725 8134 8777 8186
rect 8789 8134 8841 8186
rect 8853 8134 8905 8186
rect 6092 8032 6144 8084
rect 8024 8032 8076 8084
rect 9128 8032 9180 8084
rect 848 7828 900 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 2596 7760 2648 7812
rect 8116 7964 8168 8016
rect 8300 7964 8352 8016
rect 5724 7896 5776 7948
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 6000 7828 6052 7880
rect 6184 7760 6236 7812
rect 6276 7803 6328 7812
rect 6276 7769 6285 7803
rect 6285 7769 6319 7803
rect 6319 7769 6328 7803
rect 6276 7760 6328 7769
rect 3792 7692 3844 7744
rect 5356 7692 5408 7744
rect 5816 7735 5868 7744
rect 5816 7701 5825 7735
rect 5825 7701 5859 7735
rect 5859 7701 5868 7735
rect 5816 7692 5868 7701
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 8208 7896 8260 7948
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8392 7871 8444 7880
rect 8392 7837 8402 7871
rect 8402 7837 8444 7871
rect 8392 7828 8444 7837
rect 9036 7828 9088 7880
rect 9128 7692 9180 7744
rect 2702 7590 2754 7642
rect 2766 7590 2818 7642
rect 2830 7590 2882 7642
rect 2894 7590 2946 7642
rect 2958 7590 3010 7642
rect 4887 7590 4939 7642
rect 4951 7590 5003 7642
rect 5015 7590 5067 7642
rect 5079 7590 5131 7642
rect 5143 7590 5195 7642
rect 7072 7590 7124 7642
rect 7136 7590 7188 7642
rect 7200 7590 7252 7642
rect 7264 7590 7316 7642
rect 7328 7590 7380 7642
rect 9257 7590 9309 7642
rect 9321 7590 9373 7642
rect 9385 7590 9437 7642
rect 9449 7590 9501 7642
rect 9513 7590 9565 7642
rect 2688 7488 2740 7540
rect 3884 7488 3936 7540
rect 3976 7488 4028 7540
rect 4620 7488 4672 7540
rect 5356 7488 5408 7540
rect 2412 7420 2464 7472
rect 2412 7284 2464 7336
rect 3056 7284 3108 7336
rect 3792 7395 3844 7404
rect 3792 7361 3801 7395
rect 3801 7361 3835 7395
rect 3835 7361 3844 7395
rect 5816 7420 5868 7472
rect 8392 7420 8444 7472
rect 3792 7352 3844 7361
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 1952 7148 2004 7200
rect 4712 7284 4764 7336
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5540 7284 5592 7336
rect 4160 7216 4212 7268
rect 6920 7216 6972 7268
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 8024 7284 8076 7336
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 4804 7148 4856 7200
rect 6276 7148 6328 7200
rect 7472 7148 7524 7200
rect 8300 7284 8352 7336
rect 9220 7148 9272 7200
rect 2042 7046 2094 7098
rect 2106 7046 2158 7098
rect 2170 7046 2222 7098
rect 2234 7046 2286 7098
rect 2298 7046 2350 7098
rect 4227 7046 4279 7098
rect 4291 7046 4343 7098
rect 4355 7046 4407 7098
rect 4419 7046 4471 7098
rect 4483 7046 4535 7098
rect 6412 7046 6464 7098
rect 6476 7046 6528 7098
rect 6540 7046 6592 7098
rect 6604 7046 6656 7098
rect 6668 7046 6720 7098
rect 8597 7046 8649 7098
rect 8661 7046 8713 7098
rect 8725 7046 8777 7098
rect 8789 7046 8841 7098
rect 8853 7046 8905 7098
rect 1860 6944 1912 6996
rect 1584 6876 1636 6928
rect 2504 6876 2556 6928
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 5448 6944 5500 6996
rect 9036 6944 9088 6996
rect 2688 6808 2740 6860
rect 5356 6876 5408 6928
rect 5540 6876 5592 6928
rect 6736 6876 6788 6928
rect 1308 6672 1360 6724
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 3056 6740 3108 6792
rect 2504 6672 2556 6724
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 9220 6851 9272 6860
rect 9220 6817 9229 6851
rect 9229 6817 9263 6851
rect 9263 6817 9272 6851
rect 9220 6808 9272 6817
rect 9588 6808 9640 6860
rect 1676 6604 1728 6656
rect 1860 6604 1912 6656
rect 2136 6604 2188 6656
rect 3332 6672 3384 6724
rect 3884 6740 3936 6792
rect 4252 6740 4304 6792
rect 4896 6740 4948 6792
rect 5264 6740 5316 6792
rect 5724 6740 5776 6792
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 8116 6740 8168 6792
rect 7840 6672 7892 6724
rect 8944 6672 8996 6724
rect 3608 6604 3660 6656
rect 4620 6604 4672 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7932 6604 7984 6656
rect 8024 6604 8076 6656
rect 9128 6604 9180 6656
rect 2702 6502 2754 6554
rect 2766 6502 2818 6554
rect 2830 6502 2882 6554
rect 2894 6502 2946 6554
rect 2958 6502 3010 6554
rect 4887 6502 4939 6554
rect 4951 6502 5003 6554
rect 5015 6502 5067 6554
rect 5079 6502 5131 6554
rect 5143 6502 5195 6554
rect 7072 6502 7124 6554
rect 7136 6502 7188 6554
rect 7200 6502 7252 6554
rect 7264 6502 7316 6554
rect 7328 6502 7380 6554
rect 9257 6502 9309 6554
rect 9321 6502 9373 6554
rect 9385 6502 9437 6554
rect 9449 6502 9501 6554
rect 9513 6502 9565 6554
rect 1952 6400 2004 6452
rect 2412 6400 2464 6452
rect 1860 6375 1912 6384
rect 1860 6341 1877 6375
rect 1877 6341 1912 6375
rect 1860 6332 1912 6341
rect 5724 6332 5776 6384
rect 848 6264 900 6316
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 1768 6196 1820 6248
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 3148 6196 3200 6248
rect 4252 6196 4304 6248
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 6092 6264 6144 6316
rect 8484 6264 8536 6316
rect 5264 6128 5316 6180
rect 8116 6196 8168 6248
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 5724 6060 5776 6112
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 7472 6171 7524 6180
rect 7472 6137 7481 6171
rect 7481 6137 7515 6171
rect 7515 6137 7524 6171
rect 7472 6128 7524 6137
rect 8484 6171 8536 6180
rect 8484 6137 8493 6171
rect 8493 6137 8527 6171
rect 8527 6137 8536 6171
rect 8484 6128 8536 6137
rect 2042 5958 2094 6010
rect 2106 5958 2158 6010
rect 2170 5958 2222 6010
rect 2234 5958 2286 6010
rect 2298 5958 2350 6010
rect 4227 5958 4279 6010
rect 4291 5958 4343 6010
rect 4355 5958 4407 6010
rect 4419 5958 4471 6010
rect 4483 5958 4535 6010
rect 6412 5958 6464 6010
rect 6476 5958 6528 6010
rect 6540 5958 6592 6010
rect 6604 5958 6656 6010
rect 6668 5958 6720 6010
rect 8597 5958 8649 6010
rect 8661 5958 8713 6010
rect 8725 5958 8777 6010
rect 8789 5958 8841 6010
rect 8853 5958 8905 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 6828 5856 6880 5908
rect 8944 5856 8996 5908
rect 4252 5788 4304 5840
rect 4804 5788 4856 5840
rect 3424 5720 3476 5772
rect 7840 5788 7892 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1492 5652 1544 5704
rect 5540 5720 5592 5772
rect 4344 5584 4396 5636
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 3332 5516 3384 5568
rect 4712 5516 4764 5568
rect 6000 5652 6052 5704
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 6644 5652 6696 5704
rect 7656 5720 7708 5772
rect 5632 5627 5684 5636
rect 5632 5593 5649 5627
rect 5649 5593 5684 5627
rect 5632 5584 5684 5593
rect 5724 5516 5776 5568
rect 6276 5584 6328 5636
rect 6828 5627 6880 5636
rect 6828 5593 6837 5627
rect 6837 5593 6871 5627
rect 6871 5593 6880 5627
rect 6828 5584 6880 5593
rect 8024 5652 8076 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8208 5652 8260 5704
rect 7472 5584 7524 5636
rect 6920 5516 6972 5568
rect 8944 5516 8996 5568
rect 9220 5584 9272 5636
rect 2702 5414 2754 5466
rect 2766 5414 2818 5466
rect 2830 5414 2882 5466
rect 2894 5414 2946 5466
rect 2958 5414 3010 5466
rect 4887 5414 4939 5466
rect 4951 5414 5003 5466
rect 5015 5414 5067 5466
rect 5079 5414 5131 5466
rect 5143 5414 5195 5466
rect 7072 5414 7124 5466
rect 7136 5414 7188 5466
rect 7200 5414 7252 5466
rect 7264 5414 7316 5466
rect 7328 5414 7380 5466
rect 9257 5414 9309 5466
rect 9321 5414 9373 5466
rect 9385 5414 9437 5466
rect 9449 5414 9501 5466
rect 9513 5414 9565 5466
rect 1492 5312 1544 5364
rect 1768 5287 1820 5296
rect 1768 5253 1777 5287
rect 1777 5253 1811 5287
rect 1811 5253 1820 5287
rect 1768 5244 1820 5253
rect 3056 5312 3108 5364
rect 4804 5312 4856 5364
rect 5632 5312 5684 5364
rect 6920 5312 6972 5364
rect 2596 5244 2648 5296
rect 2780 5287 2832 5296
rect 2780 5253 2789 5287
rect 2789 5253 2823 5287
rect 2823 5253 2832 5287
rect 2780 5244 2832 5253
rect 3148 5287 3200 5296
rect 3148 5253 3157 5287
rect 3157 5253 3191 5287
rect 3191 5253 3200 5287
rect 3148 5244 3200 5253
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 5264 5287 5316 5296
rect 5264 5253 5273 5287
rect 5273 5253 5307 5287
rect 5307 5253 5316 5287
rect 5264 5244 5316 5253
rect 6276 5244 6328 5296
rect 7380 5244 7432 5296
rect 2412 5176 2464 5185
rect 4344 5176 4396 5228
rect 4712 5176 4764 5228
rect 4804 5176 4856 5228
rect 5540 5176 5592 5228
rect 6184 5176 6236 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 1860 5108 1912 5160
rect 2504 5108 2556 5160
rect 1952 5040 2004 5092
rect 4528 5040 4580 5092
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 8024 5176 8076 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 7656 5040 7708 5092
rect 8208 5083 8260 5092
rect 8208 5049 8217 5083
rect 8217 5049 8251 5083
rect 8251 5049 8260 5083
rect 8208 5040 8260 5049
rect 3332 5015 3384 5024
rect 3332 4981 3341 5015
rect 3341 4981 3375 5015
rect 3375 4981 3384 5015
rect 3332 4972 3384 4981
rect 3700 4972 3752 5024
rect 4252 4972 4304 5024
rect 4988 4972 5040 5024
rect 6368 4972 6420 5024
rect 7748 4972 7800 5024
rect 2042 4870 2094 4922
rect 2106 4870 2158 4922
rect 2170 4870 2222 4922
rect 2234 4870 2286 4922
rect 2298 4870 2350 4922
rect 4227 4870 4279 4922
rect 4291 4870 4343 4922
rect 4355 4870 4407 4922
rect 4419 4870 4471 4922
rect 4483 4870 4535 4922
rect 6412 4870 6464 4922
rect 6476 4870 6528 4922
rect 6540 4870 6592 4922
rect 6604 4870 6656 4922
rect 6668 4870 6720 4922
rect 8597 4870 8649 4922
rect 8661 4870 8713 4922
rect 8725 4870 8777 4922
rect 8789 4870 8841 4922
rect 8853 4870 8905 4922
rect 1216 4768 1268 4820
rect 1860 4768 1912 4820
rect 2780 4768 2832 4820
rect 3792 4768 3844 4820
rect 5908 4768 5960 4820
rect 8300 4768 8352 4820
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 1308 4496 1360 4548
rect 3700 4632 3752 4684
rect 3148 4564 3200 4616
rect 2412 4496 2464 4548
rect 3056 4539 3108 4548
rect 3056 4505 3065 4539
rect 3065 4505 3099 4539
rect 3099 4505 3108 4539
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4620 4632 4672 4684
rect 6184 4700 6236 4752
rect 6920 4700 6972 4752
rect 8024 4700 8076 4752
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 8300 4632 8352 4684
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 6920 4564 6972 4616
rect 3056 4496 3108 4505
rect 6644 4496 6696 4548
rect 7380 4564 7432 4616
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 7748 4496 7800 4548
rect 4620 4428 4672 4480
rect 6828 4428 6880 4480
rect 8208 4428 8260 4480
rect 9680 4496 9732 4548
rect 2702 4326 2754 4378
rect 2766 4326 2818 4378
rect 2830 4326 2882 4378
rect 2894 4326 2946 4378
rect 2958 4326 3010 4378
rect 4887 4326 4939 4378
rect 4951 4326 5003 4378
rect 5015 4326 5067 4378
rect 5079 4326 5131 4378
rect 5143 4326 5195 4378
rect 7072 4326 7124 4378
rect 7136 4326 7188 4378
rect 7200 4326 7252 4378
rect 7264 4326 7316 4378
rect 7328 4326 7380 4378
rect 9257 4326 9309 4378
rect 9321 4326 9373 4378
rect 9385 4326 9437 4378
rect 9449 4326 9501 4378
rect 9513 4326 9565 4378
rect 6184 4224 6236 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 5448 4156 5500 4208
rect 6828 4156 6880 4208
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 5264 4088 5316 4140
rect 6644 4020 6696 4072
rect 7656 4156 7708 4208
rect 8116 4156 8168 4208
rect 5632 3952 5684 4004
rect 6736 3952 6788 4004
rect 9588 4088 9640 4140
rect 7656 4020 7708 4072
rect 7932 4063 7984 4072
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 8208 4020 8260 4072
rect 8300 4063 8352 4072
rect 8300 4029 8309 4063
rect 8309 4029 8343 4063
rect 8343 4029 8352 4063
rect 8300 4020 8352 4029
rect 9680 4020 9732 4072
rect 2872 3884 2924 3936
rect 3148 3884 3200 3936
rect 4068 3884 4120 3936
rect 4896 3884 4948 3936
rect 6276 3884 6328 3936
rect 7564 3884 7616 3936
rect 8944 3884 8996 3936
rect 2042 3782 2094 3834
rect 2106 3782 2158 3834
rect 2170 3782 2222 3834
rect 2234 3782 2286 3834
rect 2298 3782 2350 3834
rect 4227 3782 4279 3834
rect 4291 3782 4343 3834
rect 4355 3782 4407 3834
rect 4419 3782 4471 3834
rect 4483 3782 4535 3834
rect 6412 3782 6464 3834
rect 6476 3782 6528 3834
rect 6540 3782 6592 3834
rect 6604 3782 6656 3834
rect 6668 3782 6720 3834
rect 8597 3782 8649 3834
rect 8661 3782 8713 3834
rect 8725 3782 8777 3834
rect 8789 3782 8841 3834
rect 8853 3782 8905 3834
rect 1584 3680 1636 3732
rect 2044 3680 2096 3732
rect 3332 3680 3384 3732
rect 4252 3680 4304 3732
rect 5356 3723 5408 3732
rect 5356 3689 5365 3723
rect 5365 3689 5399 3723
rect 5399 3689 5408 3723
rect 5356 3680 5408 3689
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 3240 3612 3292 3664
rect 6276 3680 6328 3732
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 3516 3544 3568 3596
rect 2872 3408 2924 3460
rect 3240 3476 3292 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 5724 3544 5776 3596
rect 5264 3476 5316 3528
rect 5356 3476 5408 3528
rect 6184 3476 6236 3528
rect 7564 3544 7616 3596
rect 8392 3544 8444 3596
rect 9680 3544 9732 3596
rect 1952 3340 2004 3392
rect 2596 3340 2648 3392
rect 4620 3408 4672 3460
rect 4896 3408 4948 3460
rect 3056 3340 3108 3392
rect 3332 3340 3384 3392
rect 4436 3340 4488 3392
rect 4988 3340 5040 3392
rect 7196 3408 7248 3460
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7840 3476 7892 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8300 3476 8352 3528
rect 7472 3408 7524 3460
rect 7564 3408 7616 3460
rect 9036 3408 9088 3460
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 7748 3340 7800 3392
rect 8116 3340 8168 3392
rect 2702 3238 2754 3290
rect 2766 3238 2818 3290
rect 2830 3238 2882 3290
rect 2894 3238 2946 3290
rect 2958 3238 3010 3290
rect 4887 3238 4939 3290
rect 4951 3238 5003 3290
rect 5015 3238 5067 3290
rect 5079 3238 5131 3290
rect 5143 3238 5195 3290
rect 7072 3238 7124 3290
rect 7136 3238 7188 3290
rect 7200 3238 7252 3290
rect 7264 3238 7316 3290
rect 7328 3238 7380 3290
rect 9257 3238 9309 3290
rect 9321 3238 9373 3290
rect 9385 3238 9437 3290
rect 9449 3238 9501 3290
rect 9513 3238 9565 3290
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 3332 3068 3384 3120
rect 2780 3000 2832 3052
rect 2596 2932 2648 2984
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 4620 3068 4672 3120
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 4804 3000 4856 3052
rect 5448 3136 5500 3188
rect 6092 3136 6144 3188
rect 7472 3136 7524 3188
rect 7840 3179 7892 3188
rect 7840 3145 7849 3179
rect 7849 3145 7883 3179
rect 7883 3145 7892 3179
rect 7840 3136 7892 3145
rect 7932 3136 7984 3188
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 5816 3068 5868 3120
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 7472 3000 7524 3052
rect 3516 2932 3568 2984
rect 7656 3000 7708 3052
rect 8024 2932 8076 2984
rect 8300 2975 8352 2984
rect 8300 2941 8309 2975
rect 8309 2941 8343 2975
rect 8343 2941 8352 2975
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 9036 3111 9088 3120
rect 9036 3077 9045 3111
rect 9045 3077 9079 3111
rect 9079 3077 9088 3111
rect 9036 3068 9088 3077
rect 8300 2932 8352 2941
rect 2504 2864 2556 2916
rect 4160 2864 4212 2916
rect 4252 2864 4304 2916
rect 6920 2864 6972 2916
rect 7840 2864 7892 2916
rect 6276 2796 6328 2848
rect 8576 2796 8628 2848
rect 2042 2694 2094 2746
rect 2106 2694 2158 2746
rect 2170 2694 2222 2746
rect 2234 2694 2286 2746
rect 2298 2694 2350 2746
rect 4227 2694 4279 2746
rect 4291 2694 4343 2746
rect 4355 2694 4407 2746
rect 4419 2694 4471 2746
rect 4483 2694 4535 2746
rect 6412 2694 6464 2746
rect 6476 2694 6528 2746
rect 6540 2694 6592 2746
rect 6604 2694 6656 2746
rect 6668 2694 6720 2746
rect 8597 2694 8649 2746
rect 8661 2694 8713 2746
rect 8725 2694 8777 2746
rect 8789 2694 8841 2746
rect 8853 2694 8905 2746
rect 2780 2592 2832 2644
rect 3056 2592 3108 2644
rect 3976 2592 4028 2644
rect 4804 2592 4856 2644
rect 5264 2592 5316 2644
rect 8024 2592 8076 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 8484 2592 8536 2644
rect 3240 2388 3292 2440
rect 3884 2388 3936 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5264 2388 5316 2440
rect 6276 2388 6328 2440
rect 4528 2320 4580 2372
rect 5816 2320 5868 2372
rect 6920 2252 6972 2304
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8392 2388 8444 2440
rect 7748 2252 7800 2304
rect 2702 2150 2754 2202
rect 2766 2150 2818 2202
rect 2830 2150 2882 2202
rect 2894 2150 2946 2202
rect 2958 2150 3010 2202
rect 4887 2150 4939 2202
rect 4951 2150 5003 2202
rect 5015 2150 5067 2202
rect 5079 2150 5131 2202
rect 5143 2150 5195 2202
rect 7072 2150 7124 2202
rect 7136 2150 7188 2202
rect 7200 2150 7252 2202
rect 7264 2150 7316 2202
rect 7328 2150 7380 2202
rect 9257 2150 9309 2202
rect 9321 2150 9373 2202
rect 9385 2150 9437 2202
rect 9449 2150 9501 2202
rect 9513 2150 9565 2202
<< metal2 >>
rect 3882 12308 3938 13108
rect 5170 12308 5226 13108
rect 5814 12308 5870 13108
rect 6458 12308 6514 13108
rect 7746 12308 7802 13108
rect 8390 12308 8446 13108
rect 2702 10908 3010 10917
rect 2702 10906 2708 10908
rect 2764 10906 2788 10908
rect 2844 10906 2868 10908
rect 2924 10906 2948 10908
rect 3004 10906 3010 10908
rect 2764 10854 2766 10906
rect 2946 10854 2948 10906
rect 2702 10852 2708 10854
rect 2764 10852 2788 10854
rect 2844 10852 2868 10854
rect 2924 10852 2948 10854
rect 3004 10852 3010 10854
rect 2702 10843 3010 10852
rect 3896 10826 3924 12308
rect 5184 11098 5212 12308
rect 5184 11070 5304 11098
rect 4887 10908 5195 10917
rect 4887 10906 4893 10908
rect 4949 10906 4973 10908
rect 5029 10906 5053 10908
rect 5109 10906 5133 10908
rect 5189 10906 5195 10908
rect 4949 10854 4951 10906
rect 5131 10854 5133 10906
rect 4887 10852 4893 10854
rect 4949 10852 4973 10854
rect 5029 10852 5053 10854
rect 5109 10852 5133 10854
rect 5189 10852 5195 10854
rect 4887 10843 5195 10852
rect 3424 10804 3476 10810
rect 3344 10764 3424 10792
rect 2042 10364 2350 10373
rect 2042 10362 2048 10364
rect 2104 10362 2128 10364
rect 2184 10362 2208 10364
rect 2264 10362 2288 10364
rect 2344 10362 2350 10364
rect 2104 10310 2106 10362
rect 2286 10310 2288 10362
rect 2042 10308 2048 10310
rect 2104 10308 2128 10310
rect 2184 10308 2208 10310
rect 2264 10308 2288 10310
rect 2344 10308 2350 10310
rect 2042 10299 2350 10308
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 1398 9616 1454 9625
rect 2608 9586 2636 9862
rect 2702 9820 3010 9829
rect 2702 9818 2708 9820
rect 2764 9818 2788 9820
rect 2844 9818 2868 9820
rect 2924 9818 2948 9820
rect 3004 9818 3010 9820
rect 2764 9766 2766 9818
rect 2946 9766 2948 9818
rect 2702 9764 2708 9766
rect 2764 9764 2788 9766
rect 2844 9764 2868 9766
rect 2924 9764 2948 9766
rect 3004 9764 3010 9766
rect 2702 9755 3010 9764
rect 3160 9586 3188 9862
rect 3344 9586 3372 10764
rect 3896 10798 4016 10826
rect 5276 10810 5304 11070
rect 3424 10746 3476 10752
rect 3988 10742 4016 10798
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 9722 3464 10406
rect 3620 10130 3648 10542
rect 3712 10130 3740 10678
rect 5828 10674 5856 12308
rect 6472 10690 6500 12308
rect 7072 10908 7380 10917
rect 7072 10906 7078 10908
rect 7134 10906 7158 10908
rect 7214 10906 7238 10908
rect 7294 10906 7318 10908
rect 7374 10906 7380 10908
rect 7134 10854 7136 10906
rect 7316 10854 7318 10906
rect 7072 10852 7078 10854
rect 7134 10852 7158 10854
rect 7214 10852 7238 10854
rect 7294 10852 7318 10854
rect 7374 10852 7380 10854
rect 7072 10843 7380 10852
rect 7760 10742 7788 12308
rect 7748 10736 7800 10742
rect 6472 10674 6592 10690
rect 7748 10678 7800 10684
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 6092 10668 6144 10674
rect 6472 10668 6604 10674
rect 6472 10662 6552 10668
rect 6092 10610 6144 10616
rect 6552 10610 6604 10616
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3988 10062 4016 10406
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 4080 9586 4108 10610
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 4227 10364 4535 10373
rect 4227 10362 4233 10364
rect 4289 10362 4313 10364
rect 4369 10362 4393 10364
rect 4449 10362 4473 10364
rect 4529 10362 4535 10364
rect 4289 10310 4291 10362
rect 4471 10310 4473 10362
rect 4227 10308 4233 10310
rect 4289 10308 4313 10310
rect 4369 10308 4393 10310
rect 4449 10308 4473 10310
rect 4529 10308 4535 10310
rect 4227 10299 4535 10308
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 1398 9551 1454 9560
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2780 9580 2832 9586
rect 3148 9580 3200 9586
rect 2832 9540 3096 9568
rect 2780 9522 2832 9528
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2042 9276 2350 9285
rect 2042 9274 2048 9276
rect 2104 9274 2128 9276
rect 2184 9274 2208 9276
rect 2264 9274 2288 9276
rect 2344 9274 2350 9276
rect 2104 9222 2106 9274
rect 2286 9222 2288 9274
rect 2042 9220 2048 9222
rect 2104 9220 2128 9222
rect 2184 9220 2208 9222
rect 2264 9220 2288 9222
rect 2344 9220 2350 9222
rect 2042 9211 2350 9220
rect 2424 9110 2452 9318
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 2412 9104 2464 9110
rect 900 9072 902 9081
rect 2412 9046 2464 9052
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 846 9007 902 9016
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1780 8634 1808 8910
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1320 6730 1348 8434
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1872 7002 1900 8978
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2516 8498 2544 9046
rect 2608 9042 2636 9522
rect 3068 9382 3096 9540
rect 3148 9522 3200 9528
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2976 8906 3004 9318
rect 3344 8906 3372 9522
rect 4172 9330 4200 9998
rect 4540 9586 4568 10066
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4080 9302 4200 9330
rect 4080 9194 4108 9302
rect 4227 9276 4535 9285
rect 4227 9274 4233 9276
rect 4289 9274 4313 9276
rect 4369 9274 4393 9276
rect 4449 9274 4473 9276
rect 4529 9274 4535 9276
rect 4289 9222 4291 9274
rect 4471 9222 4473 9274
rect 4227 9220 4233 9222
rect 4289 9220 4313 9222
rect 4369 9220 4393 9222
rect 4449 9220 4473 9222
rect 4529 9220 4535 9222
rect 4227 9211 4535 9220
rect 4080 9166 4200 9194
rect 4632 9178 4660 10542
rect 5276 10198 5304 10542
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4816 9654 4844 9998
rect 4887 9820 5195 9829
rect 4887 9818 4893 9820
rect 4949 9818 4973 9820
rect 5029 9818 5053 9820
rect 5109 9818 5133 9820
rect 5189 9818 5195 9820
rect 4949 9766 4951 9818
rect 5131 9766 5133 9818
rect 4887 9764 4893 9766
rect 4949 9764 4973 9766
rect 5029 9764 5053 9766
rect 5109 9764 5133 9766
rect 5189 9764 5195 9766
rect 4887 9755 5195 9764
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 2702 8732 3010 8741
rect 2702 8730 2708 8732
rect 2764 8730 2788 8732
rect 2844 8730 2868 8732
rect 2924 8730 2948 8732
rect 3004 8730 3010 8732
rect 2764 8678 2766 8730
rect 2946 8678 2948 8730
rect 2702 8676 2708 8678
rect 2764 8676 2788 8678
rect 2844 8676 2868 8678
rect 2924 8676 2948 8678
rect 3004 8676 3010 8678
rect 2702 8667 3010 8676
rect 3804 8498 3832 8774
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 2042 8188 2350 8197
rect 2042 8186 2048 8188
rect 2104 8186 2128 8188
rect 2184 8186 2208 8188
rect 2264 8186 2288 8188
rect 2344 8186 2350 8188
rect 2104 8134 2106 8186
rect 2286 8134 2288 8186
rect 2042 8132 2048 8134
rect 2104 8132 2128 8134
rect 2184 8132 2208 8134
rect 2264 8132 2288 8134
rect 2344 8132 2350 8134
rect 2042 8123 2350 8132
rect 2608 7818 2636 8366
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2412 7472 2464 7478
rect 2464 7432 2544 7460
rect 2412 7414 2464 7420
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1584 6928 1636 6934
rect 1490 6896 1546 6905
rect 1584 6870 1636 6876
rect 1490 6831 1546 6840
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1214 4856 1270 4865
rect 1214 4791 1216 4800
rect 1268 4791 1270 4800
rect 1216 4762 1268 4768
rect 1320 4554 1348 6666
rect 1596 5914 1624 6870
rect 1872 6746 1900 6938
rect 1780 6718 1900 6746
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6322 1716 6598
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1780 6254 1808 6718
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6390 1900 6598
rect 1964 6458 1992 7142
rect 2042 7100 2350 7109
rect 2042 7098 2048 7100
rect 2104 7098 2128 7100
rect 2184 7098 2208 7100
rect 2264 7098 2288 7100
rect 2344 7098 2350 7100
rect 2104 7046 2106 7098
rect 2286 7046 2288 7098
rect 2042 7044 2048 7046
rect 2104 7044 2128 7046
rect 2184 7044 2208 7046
rect 2264 7044 2288 7046
rect 2344 7044 2350 7046
rect 2042 7035 2350 7044
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 2148 6322 2176 6598
rect 2424 6458 2452 7278
rect 2516 6934 2544 7432
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2608 6798 2636 7754
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 2702 7644 3010 7653
rect 2702 7642 2708 7644
rect 2764 7642 2788 7644
rect 2844 7642 2868 7644
rect 2924 7642 2948 7644
rect 3004 7642 3010 7644
rect 2764 7590 2766 7642
rect 2946 7590 2948 7642
rect 2702 7588 2708 7590
rect 2764 7588 2788 7590
rect 2844 7588 2868 7590
rect 2924 7588 2948 7590
rect 3004 7588 3010 7590
rect 2702 7579 3010 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2700 6866 2728 7482
rect 3804 7410 3832 7686
rect 3988 7546 4016 8366
rect 4172 8242 4200 9166
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4724 8498 4752 9318
rect 4816 8974 4844 9590
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 9110 4936 9318
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8566 4844 8910
rect 5092 8838 5120 9386
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4887 8732 5195 8741
rect 4887 8730 4893 8732
rect 4949 8730 4973 8732
rect 5029 8730 5053 8732
rect 5109 8730 5133 8732
rect 5189 8730 5195 8732
rect 4949 8678 4951 8730
rect 5131 8678 5133 8730
rect 4887 8676 4893 8678
rect 4949 8676 4973 8678
rect 5029 8676 5053 8678
rect 5109 8676 5133 8678
rect 5189 8676 5195 8678
rect 4887 8667 5195 8676
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4080 8214 4200 8242
rect 4080 8106 4108 8214
rect 4227 8188 4535 8197
rect 4227 8186 4233 8188
rect 4289 8186 4313 8188
rect 4369 8186 4393 8188
rect 4449 8186 4473 8188
rect 4529 8186 4535 8188
rect 4289 8134 4291 8186
rect 4471 8134 4473 8186
rect 4227 8132 4233 8134
rect 4289 8132 4313 8134
rect 4369 8132 4393 8134
rect 4449 8132 4473 8134
rect 4529 8132 4535 8134
rect 4227 8123 4535 8132
rect 4080 8078 4200 8106
rect 4172 7970 4200 8078
rect 4172 7942 4292 7970
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 3068 6798 3096 7278
rect 3804 6882 3832 7346
rect 3896 7002 3924 7482
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 7154 4200 7210
rect 4264 7206 4292 7942
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4632 7546 4660 7822
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4816 7460 4844 8366
rect 5092 7886 5120 8366
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7886 5212 8230
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5276 7834 5304 10134
rect 5368 10130 5396 10542
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 9586 5396 10066
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8498 5488 9318
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5460 8294 5488 8434
rect 5552 8430 5580 9454
rect 5828 9042 5856 10406
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9586 6040 9998
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5276 7806 5488 7834
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 4887 7644 5195 7653
rect 4887 7642 4893 7644
rect 4949 7642 4973 7644
rect 5029 7642 5053 7644
rect 5109 7642 5133 7644
rect 5189 7642 5195 7644
rect 4949 7590 4951 7642
rect 5131 7590 5133 7642
rect 4887 7588 4893 7590
rect 4949 7588 4973 7590
rect 5029 7588 5053 7590
rect 5109 7588 5133 7590
rect 5189 7588 5195 7590
rect 4887 7579 5195 7588
rect 5368 7546 5396 7686
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 4816 7432 4936 7460
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4080 7126 4200 7154
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4080 7018 4108 7126
rect 4227 7100 4535 7109
rect 4227 7098 4233 7100
rect 4289 7098 4313 7100
rect 4369 7098 4393 7100
rect 4449 7098 4473 7100
rect 4529 7098 4535 7100
rect 4289 7046 4291 7098
rect 4471 7046 4473 7098
rect 4227 7044 4233 7046
rect 4289 7044 4313 7046
rect 4369 7044 4393 7046
rect 4449 7044 4473 7046
rect 4529 7044 4535 7046
rect 4227 7035 4535 7044
rect 3884 6996 3936 7002
rect 4080 6990 4200 7018
rect 3884 6938 3936 6944
rect 3804 6854 3924 6882
rect 3896 6798 3924 6854
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1504 5370 1532 5646
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1308 4548 1360 4554
rect 1308 4490 1360 4496
rect 1398 4176 1454 4185
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 1400 4082 1452 4088
rect 1596 3738 1624 5170
rect 1688 4622 1716 5510
rect 1780 5302 1808 6190
rect 2042 6012 2350 6021
rect 2042 6010 2048 6012
rect 2104 6010 2128 6012
rect 2184 6010 2208 6012
rect 2264 6010 2288 6012
rect 2344 6010 2350 6012
rect 2104 5958 2106 6010
rect 2286 5958 2288 6010
rect 2042 5956 2048 5958
rect 2104 5956 2128 5958
rect 2184 5956 2208 5958
rect 2264 5956 2288 5958
rect 2344 5956 2350 5958
rect 2042 5947 2350 5956
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1872 4826 1900 5102
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1964 3398 1992 5034
rect 2042 4924 2350 4933
rect 2042 4922 2048 4924
rect 2104 4922 2128 4924
rect 2184 4922 2208 4924
rect 2264 4922 2288 4924
rect 2344 4922 2350 4924
rect 2104 4870 2106 4922
rect 2286 4870 2288 4922
rect 2042 4868 2048 4870
rect 2104 4868 2128 4870
rect 2184 4868 2208 4870
rect 2264 4868 2288 4870
rect 2344 4868 2350 4870
rect 2042 4859 2350 4868
rect 2424 4554 2452 5170
rect 2516 5166 2544 6666
rect 2608 5302 2636 6734
rect 2702 6556 3010 6565
rect 2702 6554 2708 6556
rect 2764 6554 2788 6556
rect 2844 6554 2868 6556
rect 2924 6554 2948 6556
rect 3004 6554 3010 6556
rect 2764 6502 2766 6554
rect 2946 6502 2948 6554
rect 2702 6500 2708 6502
rect 2764 6500 2788 6502
rect 2844 6500 2868 6502
rect 2924 6500 2948 6502
rect 3004 6500 3010 6502
rect 2702 6491 3010 6500
rect 2702 5468 3010 5477
rect 2702 5466 2708 5468
rect 2764 5466 2788 5468
rect 2844 5466 2868 5468
rect 2924 5466 2948 5468
rect 3004 5466 3010 5468
rect 2764 5414 2766 5466
rect 2946 5414 2948 5466
rect 2702 5412 2708 5414
rect 2764 5412 2788 5414
rect 2844 5412 2868 5414
rect 2924 5412 2948 5414
rect 3004 5412 3010 5414
rect 2702 5403 3010 5412
rect 3068 5370 3096 6734
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 6322 3372 6666
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6322 3648 6598
rect 4172 6322 4200 6990
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4264 6254 4292 6734
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3160 5302 3188 6190
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5778 3464 6054
rect 4227 6012 4535 6021
rect 4227 6010 4233 6012
rect 4289 6010 4313 6012
rect 4369 6010 4393 6012
rect 4449 6010 4473 6012
rect 4529 6010 4535 6012
rect 4289 5958 4291 6010
rect 4471 5958 4473 6010
rect 4227 5956 4233 5958
rect 4289 5956 4313 5958
rect 4369 5956 4393 5958
rect 4449 5956 4473 5958
rect 4529 5956 4535 5958
rect 4227 5947 4535 5956
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 2596 5296 2648 5302
rect 2594 5264 2596 5273
rect 2780 5296 2832 5302
rect 2648 5264 2650 5273
rect 2780 5238 2832 5244
rect 3148 5296 3200 5302
rect 3200 5256 3280 5284
rect 3148 5238 3200 5244
rect 2594 5199 2650 5208
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2792 4826 2820 5238
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2702 4380 3010 4389
rect 2702 4378 2708 4380
rect 2764 4378 2788 4380
rect 2844 4378 2868 4380
rect 2924 4378 2948 4380
rect 3004 4378 3010 4380
rect 2764 4326 2766 4378
rect 2946 4326 2948 4378
rect 2702 4324 2708 4326
rect 2764 4324 2788 4326
rect 2844 4324 2868 4326
rect 2924 4324 2948 4326
rect 3004 4324 3010 4326
rect 2702 4315 3010 4324
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2042 3836 2350 3845
rect 2042 3834 2048 3836
rect 2104 3834 2128 3836
rect 2184 3834 2208 3836
rect 2264 3834 2288 3836
rect 2344 3834 2350 3836
rect 2104 3782 2106 3834
rect 2286 3782 2288 3834
rect 2042 3780 2048 3782
rect 2104 3780 2128 3782
rect 2184 3780 2208 3782
rect 2264 3780 2288 3782
rect 2344 3780 2350 3782
rect 2042 3771 2350 3780
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2056 3534 2084 3674
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2516 2922 2544 3470
rect 2884 3466 2912 3878
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 3068 3398 3096 4490
rect 3160 3942 3188 4558
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2608 2990 2636 3334
rect 2702 3292 3010 3301
rect 2702 3290 2708 3292
rect 2764 3290 2788 3292
rect 2844 3290 2868 3292
rect 2924 3290 2948 3292
rect 3004 3290 3010 3292
rect 2764 3238 2766 3290
rect 2946 3238 2948 3290
rect 2702 3236 2708 3238
rect 2764 3236 2788 3238
rect 2844 3236 2868 3238
rect 2924 3236 2948 3238
rect 3004 3236 3010 3238
rect 2702 3227 3010 3236
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2042 2748 2350 2757
rect 2042 2746 2048 2748
rect 2104 2746 2128 2748
rect 2184 2746 2208 2748
rect 2264 2746 2288 2748
rect 2344 2746 2350 2748
rect 2104 2694 2106 2746
rect 2286 2694 2288 2746
rect 2042 2692 2048 2694
rect 2104 2692 2128 2694
rect 2184 2692 2208 2694
rect 2264 2692 2288 2694
rect 2344 2692 2350 2694
rect 2042 2683 2350 2692
rect 2792 2650 2820 2994
rect 3068 2650 3096 3334
rect 3160 3058 3188 3878
rect 3252 3670 3280 5256
rect 3344 5030 3372 5510
rect 4264 5030 4292 5782
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4356 5234 4384 5578
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4526 5128 4582 5137
rect 4526 5063 4528 5072
rect 4580 5063 4582 5072
rect 4528 5034 4580 5040
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3344 3738 3372 4966
rect 3712 4690 3740 4966
rect 4227 4924 4535 4933
rect 4227 4922 4233 4924
rect 4289 4922 4313 4924
rect 4369 4922 4393 4924
rect 4449 4922 4473 4924
rect 4529 4922 4535 4924
rect 4289 4870 4291 4922
rect 4471 4870 4473 4922
rect 4227 4868 4233 4870
rect 4289 4868 4313 4870
rect 4369 4868 4393 4870
rect 4449 4868 4473 4870
rect 4529 4868 4535 4870
rect 4227 4859 4535 4868
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3804 4622 3832 4762
rect 4632 4690 4660 6598
rect 4724 5574 4752 7278
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 5846 4844 7142
rect 4908 6798 4936 7432
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5368 6934 5396 7346
rect 5460 7002 5488 7806
rect 5552 7342 5580 8230
rect 5644 7410 5672 8230
rect 5736 7954 5764 8910
rect 5828 8498 5856 8978
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6012 7886 6040 8298
rect 6104 8090 6132 10610
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 9586 6224 10406
rect 6412 10364 6720 10373
rect 6412 10362 6418 10364
rect 6474 10362 6498 10364
rect 6554 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6720 10364
rect 6474 10310 6476 10362
rect 6656 10310 6658 10362
rect 6412 10308 6418 10310
rect 6474 10308 6498 10310
rect 6554 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6720 10310
rect 6412 10299 6720 10308
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9994 6776 10066
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9654 6316 9862
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6748 9586 6776 9930
rect 6932 9586 6960 10474
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10062 7052 10406
rect 7944 10130 7972 10542
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7072 9820 7380 9829
rect 7072 9818 7078 9820
rect 7134 9818 7158 9820
rect 7214 9818 7238 9820
rect 7294 9818 7318 9820
rect 7374 9818 7380 9820
rect 7134 9766 7136 9818
rect 7316 9766 7318 9818
rect 7072 9764 7078 9766
rect 7134 9764 7158 9766
rect 7214 9764 7238 9766
rect 7294 9764 7318 9766
rect 7374 9764 7380 9766
rect 7072 9755 7380 9764
rect 7484 9586 7512 9998
rect 7760 9722 7788 9998
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 6196 8430 6224 9386
rect 6412 9276 6720 9285
rect 6412 9274 6418 9276
rect 6474 9274 6498 9276
rect 6554 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6720 9276
rect 6474 9222 6476 9274
rect 6656 9222 6658 9274
rect 6412 9220 6418 9222
rect 6474 9220 6498 9222
rect 6554 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6720 9222
rect 6412 9211 6720 9220
rect 6840 8566 6868 9386
rect 7072 8732 7380 8741
rect 7072 8730 7078 8732
rect 7134 8730 7158 8732
rect 7214 8730 7238 8732
rect 7294 8730 7318 8732
rect 7374 8730 7380 8732
rect 7134 8678 7136 8730
rect 7316 8678 7318 8730
rect 7072 8676 7078 8678
rect 7134 8676 7158 8678
rect 7214 8676 7238 8678
rect 7294 8676 7318 8678
rect 7374 8676 7380 8678
rect 7072 8667 7380 8676
rect 7484 8634 7512 9386
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 7102 8528 7158 8537
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6552 8492 6604 8498
rect 7012 8492 7064 8498
rect 6552 8434 6604 8440
rect 6932 8452 7012 8480
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 7478 5856 7686
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4887 6556 5195 6565
rect 4887 6554 4893 6556
rect 4949 6554 4973 6556
rect 5029 6554 5053 6556
rect 5109 6554 5133 6556
rect 5189 6554 5195 6556
rect 4949 6502 4951 6554
rect 5131 6502 5133 6554
rect 4887 6500 4893 6502
rect 4949 6500 4973 6502
rect 5029 6500 5053 6502
rect 5109 6500 5133 6502
rect 5189 6500 5195 6502
rect 4887 6491 5195 6500
rect 5276 6186 5304 6734
rect 5552 6322 5580 6870
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6390 5764 6734
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 5552 5778 5580 6258
rect 5736 6118 5764 6326
rect 6012 6118 6040 7822
rect 6196 7818 6224 8366
rect 6288 7818 6316 8434
rect 6564 8294 6592 8434
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6412 8188 6720 8197
rect 6412 8186 6418 8188
rect 6474 8186 6498 8188
rect 6554 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6720 8188
rect 6474 8134 6476 8186
rect 6656 8134 6658 8186
rect 6412 8132 6418 8134
rect 6474 8132 6498 8134
rect 6554 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6720 8134
rect 6412 8123 6720 8132
rect 6932 7886 6960 8452
rect 7102 8463 7158 8472
rect 7380 8492 7432 8498
rect 7012 8434 7064 8440
rect 7116 8362 7144 8463
rect 7380 8434 7432 8440
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7392 7993 7420 8434
rect 7378 7984 7434 7993
rect 7378 7919 7434 7928
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6288 7206 6316 7754
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6610 6316 7142
rect 6412 7100 6720 7109
rect 6412 7098 6418 7100
rect 6474 7098 6498 7100
rect 6554 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6720 7100
rect 6474 7046 6476 7098
rect 6656 7046 6658 7098
rect 6412 7044 6418 7046
rect 6474 7044 6498 7046
rect 6554 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6720 7046
rect 6412 7035 6720 7044
rect 6748 6934 6776 7822
rect 6932 7274 6960 7822
rect 7072 7644 7380 7653
rect 7072 7642 7078 7644
rect 7134 7642 7158 7644
rect 7214 7642 7238 7644
rect 7294 7642 7318 7644
rect 7374 7642 7380 7644
rect 7134 7590 7136 7642
rect 7316 7590 7318 7642
rect 7072 7588 7078 7590
rect 7134 7588 7158 7590
rect 7214 7588 7238 7590
rect 7294 7588 7318 7590
rect 7374 7588 7380 7590
rect 7072 7579 7380 7588
rect 7378 7440 7434 7449
rect 7378 7375 7434 7384
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 7392 6662 7420 7375
rect 7484 7206 7512 8570
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7576 6798 7604 9046
rect 7668 7993 7696 9454
rect 7760 9382 7788 9522
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7654 7984 7710 7993
rect 7654 7919 7710 7928
rect 7748 7880 7800 7886
rect 7852 7868 7880 8910
rect 7800 7840 7880 7868
rect 7748 7822 7800 7828
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 6196 6582 6316 6610
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4887 5468 5195 5477
rect 4887 5466 4893 5468
rect 4949 5466 4973 5468
rect 5029 5466 5053 5468
rect 5109 5466 5133 5468
rect 5189 5466 5195 5468
rect 4949 5414 4951 5466
rect 5131 5414 5133 5466
rect 4887 5412 4893 5414
rect 4949 5412 4973 5414
rect 5029 5412 5053 5414
rect 5109 5412 5133 5414
rect 5189 5412 5195 5414
rect 4887 5403 5195 5412
rect 4804 5364 4856 5370
rect 4724 5324 4804 5352
rect 4724 5234 4752 5324
rect 4804 5306 4856 5312
rect 5264 5296 5316 5302
rect 5262 5264 5264 5273
rect 5316 5264 5318 5273
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4804 5228 4856 5234
rect 5552 5234 5580 5714
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5370 5672 5578
rect 5736 5574 5764 6054
rect 6012 5710 6040 6054
rect 6104 5914 6132 6258
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5262 5199 5318 5208
rect 5540 5228 5592 5234
rect 4804 5170 4856 5176
rect 5540 5170 5592 5176
rect 4710 5128 4766 5137
rect 4710 5063 4766 5072
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3252 3194 3280 3470
rect 3344 3398 3372 3674
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3344 3126 3372 3334
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3528 2990 3556 3538
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3988 2650 4016 3470
rect 4080 2904 4108 3878
rect 4227 3836 4535 3845
rect 4227 3834 4233 3836
rect 4289 3834 4313 3836
rect 4369 3834 4393 3836
rect 4449 3834 4473 3836
rect 4529 3834 4535 3836
rect 4289 3782 4291 3834
rect 4471 3782 4473 3834
rect 4227 3780 4233 3782
rect 4289 3780 4313 3782
rect 4369 3780 4393 3782
rect 4449 3780 4473 3782
rect 4529 3780 4535 3782
rect 4227 3771 4535 3780
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4264 3194 4292 3674
rect 4632 3466 4660 4422
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4264 2922 4292 3130
rect 4448 3058 4476 3334
rect 4632 3126 4660 3402
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4160 2916 4212 2922
rect 4080 2876 4160 2904
rect 4160 2858 4212 2864
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4227 2748 4535 2757
rect 4227 2746 4233 2748
rect 4289 2746 4313 2748
rect 4369 2746 4393 2748
rect 4449 2746 4473 2748
rect 4529 2746 4535 2748
rect 4289 2694 4291 2746
rect 4471 2694 4473 2746
rect 4227 2692 4233 2694
rect 4289 2692 4313 2694
rect 4369 2692 4393 2694
rect 4449 2692 4473 2694
rect 4529 2692 4535 2694
rect 4227 2683 4535 2692
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4724 2446 4752 5063
rect 4816 4622 4844 5170
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 4622 5028 4966
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4816 4162 4844 4558
rect 4887 4380 5195 4389
rect 4887 4378 4893 4380
rect 4949 4378 4973 4380
rect 5029 4378 5053 4380
rect 5109 4378 5133 4380
rect 5189 4378 5195 4380
rect 4949 4326 4951 4378
rect 5131 4326 5133 4378
rect 4887 4324 4893 4326
rect 4949 4324 4973 4326
rect 5029 4324 5053 4326
rect 5109 4324 5133 4326
rect 5189 4324 5195 4326
rect 4887 4315 5195 4324
rect 4816 4134 4936 4162
rect 4908 3942 4936 4134
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3466 4936 3878
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 5000 3398 5028 4082
rect 5276 3534 5304 4082
rect 5368 3738 5396 5102
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5368 3534 5396 3674
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4887 3292 5195 3301
rect 4887 3290 4893 3292
rect 4949 3290 4973 3292
rect 5029 3290 5053 3292
rect 5109 3290 5133 3292
rect 5189 3290 5195 3292
rect 4949 3238 4951 3290
rect 5131 3238 5133 3290
rect 4887 3236 4893 3238
rect 4949 3236 4973 3238
rect 5029 3236 5053 3238
rect 5109 3236 5133 3238
rect 5189 3236 5195 3238
rect 4887 3227 5195 3236
rect 5276 3058 5304 3470
rect 5460 3194 5488 4150
rect 5644 4010 5672 5102
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5736 3602 5764 5510
rect 6196 5234 6224 6582
rect 7072 6556 7380 6565
rect 7072 6554 7078 6556
rect 7134 6554 7158 6556
rect 7214 6554 7238 6556
rect 7294 6554 7318 6556
rect 7374 6554 7380 6556
rect 7134 6502 7136 6554
rect 7316 6502 7318 6554
rect 7072 6500 7078 6502
rect 7134 6500 7158 6502
rect 7214 6500 7238 6502
rect 7294 6500 7318 6502
rect 7374 6500 7380 6502
rect 7072 6491 7380 6500
rect 7470 6216 7526 6225
rect 7470 6151 7472 6160
rect 7524 6151 7526 6160
rect 7472 6122 7524 6128
rect 6412 6012 6720 6021
rect 6412 6010 6418 6012
rect 6474 6010 6498 6012
rect 6554 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6720 6012
rect 6474 5958 6476 6010
rect 6656 5958 6658 6010
rect 6412 5956 6418 5958
rect 6474 5956 6498 5958
rect 6554 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6720 5958
rect 6412 5947 6720 5956
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6288 5302 6316 5578
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5828 3126 5856 5102
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6196 4758 6224 5170
rect 6380 5030 6408 5646
rect 6656 5216 6684 5646
rect 6840 5642 6868 5850
rect 7852 5846 7880 6666
rect 7944 6662 7972 10066
rect 8128 9654 8156 10474
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 9674 8340 10406
rect 8404 10130 8432 12308
rect 9257 10908 9565 10917
rect 9257 10906 9263 10908
rect 9319 10906 9343 10908
rect 9399 10906 9423 10908
rect 9479 10906 9503 10908
rect 9559 10906 9565 10908
rect 9319 10854 9321 10906
rect 9501 10854 9503 10906
rect 9257 10852 9263 10854
rect 9319 10852 9343 10854
rect 9399 10852 9423 10854
rect 9479 10852 9503 10854
rect 9559 10852 9565 10854
rect 9257 10843 9565 10852
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8496 10062 8524 10610
rect 8597 10364 8905 10373
rect 8597 10362 8603 10364
rect 8659 10362 8683 10364
rect 8739 10362 8763 10364
rect 8819 10362 8843 10364
rect 8899 10362 8905 10364
rect 8659 10310 8661 10362
rect 8841 10310 8843 10362
rect 8597 10308 8603 10310
rect 8659 10308 8683 10310
rect 8739 10308 8763 10310
rect 8819 10308 8843 10310
rect 8899 10308 8905 10310
rect 8597 10299 8905 10308
rect 9140 10266 9168 10610
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8404 9722 8432 9930
rect 8496 9722 8524 9998
rect 9140 9994 9168 10202
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8220 9646 8340 9674
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9489 8064 9522
rect 8022 9480 8078 9489
rect 8220 9450 8248 9646
rect 8680 9586 8708 9862
rect 9140 9654 9168 9930
rect 9257 9820 9565 9829
rect 9257 9818 9263 9820
rect 9319 9818 9343 9820
rect 9399 9818 9423 9820
rect 9479 9818 9503 9820
rect 9559 9818 9565 9820
rect 9319 9766 9321 9818
rect 9501 9766 9503 9818
rect 9257 9764 9263 9766
rect 9319 9764 9343 9766
rect 9399 9764 9423 9766
rect 9479 9764 9503 9766
rect 9559 9764 9565 9766
rect 9257 9755 9565 9764
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8668 9580 8720 9586
rect 8496 9540 8668 9568
rect 8022 9415 8024 9424
rect 8076 9415 8078 9424
rect 8208 9444 8260 9450
rect 8024 9386 8076 9392
rect 8208 9386 8260 9392
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8090 8064 8774
rect 8128 8634 8156 9318
rect 8220 9042 8248 9386
rect 8496 9160 8524 9540
rect 8668 9522 8720 9528
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 8760 9512 8812 9518
rect 8758 9480 8760 9489
rect 8812 9480 8814 9489
rect 8758 9415 8814 9424
rect 8597 9276 8905 9285
rect 8597 9274 8603 9276
rect 8659 9274 8683 9276
rect 8739 9274 8763 9276
rect 8819 9274 8843 9276
rect 8899 9274 8905 9276
rect 8659 9222 8661 9274
rect 8841 9222 8843 9274
rect 8597 9220 8603 9222
rect 8659 9220 8683 9222
rect 8739 9220 8763 9222
rect 8819 9220 8843 9222
rect 8899 9220 8905 9222
rect 8597 9211 8905 9220
rect 8496 9132 8616 9160
rect 8588 9042 8616 9132
rect 9324 9042 9352 9522
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 8208 9036 8260 9042
rect 8576 9036 8628 9042
rect 8260 8996 8340 9024
rect 8208 8978 8260 8984
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8128 8022 8156 8434
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8220 7954 8248 8774
rect 8312 8566 8340 8996
rect 8576 8978 8628 8984
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9036 8968 9088 8974
rect 9220 8968 9272 8974
rect 9036 8910 9088 8916
rect 9140 8916 9220 8922
rect 9140 8910 9272 8916
rect 8404 8566 8432 8910
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 8022 8340 8298
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8404 7886 8432 8502
rect 8496 8362 8524 8910
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8588 8537 8616 8570
rect 8574 8528 8630 8537
rect 8574 8463 8630 8472
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8597 8188 8905 8197
rect 8597 8186 8603 8188
rect 8659 8186 8683 8188
rect 8739 8186 8763 8188
rect 8819 8186 8843 8188
rect 8899 8186 8905 8188
rect 8659 8134 8661 8186
rect 8841 8134 8843 8186
rect 8597 8132 8603 8134
rect 8659 8132 8683 8134
rect 8739 8132 8763 8134
rect 8819 8132 8843 8134
rect 8899 8132 8905 8134
rect 8597 8123 8905 8132
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7478 8432 7822
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8036 6662 8064 7278
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8128 6254 8156 6734
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5370 6960 5510
rect 7072 5468 7380 5477
rect 7072 5466 7078 5468
rect 7134 5466 7158 5468
rect 7214 5466 7238 5468
rect 7294 5466 7318 5468
rect 7374 5466 7380 5468
rect 7134 5414 7136 5466
rect 7316 5414 7318 5466
rect 7072 5412 7078 5414
rect 7134 5412 7158 5414
rect 7214 5412 7238 5414
rect 7294 5412 7318 5414
rect 7374 5412 7380 5414
rect 7072 5403 7380 5412
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7380 5296 7432 5302
rect 7194 5264 7250 5273
rect 6736 5228 6788 5234
rect 6656 5188 6736 5216
rect 7380 5238 7432 5244
rect 7194 5199 7196 5208
rect 6736 5170 6788 5176
rect 7248 5199 7250 5208
rect 7196 5170 7248 5176
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6412 4924 6720 4933
rect 6412 4922 6418 4924
rect 6474 4922 6498 4924
rect 6554 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6720 4924
rect 6474 4870 6476 4922
rect 6656 4870 6658 4922
rect 6412 4868 6418 4870
rect 6474 4868 6498 4870
rect 6554 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6720 4870
rect 6412 4859 6720 4868
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6196 4282 6224 4694
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6656 4078 6684 4490
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6748 4010 6776 5170
rect 6920 4752 6972 4758
rect 6840 4700 6920 4706
rect 6840 4694 6972 4700
rect 6840 4678 6960 4694
rect 6840 4622 6868 4678
rect 7392 4622 7420 5238
rect 7484 5234 7512 5578
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7668 5098 7696 5714
rect 8128 5710 8156 6190
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8036 5234 8064 5646
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7668 4622 7696 5034
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4214 6868 4422
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6288 3738 6316 3878
rect 6412 3836 6720 3845
rect 6412 3834 6418 3836
rect 6474 3834 6498 3836
rect 6554 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6720 3836
rect 6474 3782 6476 3834
rect 6656 3782 6658 3834
rect 6412 3780 6418 3782
rect 6474 3780 6498 3782
rect 6554 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6720 3782
rect 6412 3771 6720 3780
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6104 3194 6132 3334
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6196 3058 6224 3470
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 4816 2650 4844 2994
rect 5276 2650 5304 2994
rect 6932 2922 6960 4558
rect 7072 4380 7380 4389
rect 7072 4378 7078 4380
rect 7134 4378 7158 4380
rect 7214 4378 7238 4380
rect 7294 4378 7318 4380
rect 7374 4378 7380 4380
rect 7134 4326 7136 4378
rect 7316 4326 7318 4378
rect 7072 4324 7078 4326
rect 7134 4324 7158 4326
rect 7214 4324 7238 4326
rect 7294 4324 7318 4326
rect 7374 4324 7380 4326
rect 7072 4315 7380 4324
rect 7668 4214 7696 4558
rect 7760 4554 7788 4966
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 8036 4078 8064 4694
rect 8128 4214 8156 5646
rect 8220 5098 8248 5646
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8220 4622 8248 5034
rect 8312 4826 8340 7278
rect 8597 7100 8905 7109
rect 8597 7098 8603 7100
rect 8659 7098 8683 7100
rect 8739 7098 8763 7100
rect 8819 7098 8843 7100
rect 8899 7098 8905 7100
rect 8659 7046 8661 7098
rect 8841 7046 8843 7098
rect 8597 7044 8603 7046
rect 8659 7044 8683 7046
rect 8739 7044 8763 7046
rect 8819 7044 8843 7046
rect 8899 7044 8905 7046
rect 8597 7035 8905 7044
rect 8956 6866 8984 8910
rect 9048 8294 9076 8910
rect 9140 8894 9260 8910
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9140 8090 9168 8894
rect 9257 8732 9565 8741
rect 9257 8730 9263 8732
rect 9319 8730 9343 8732
rect 9399 8730 9423 8732
rect 9479 8730 9503 8732
rect 9559 8730 9565 8732
rect 9319 8678 9321 8730
rect 9501 8678 9503 8730
rect 9257 8676 9263 8678
rect 9319 8676 9343 8678
rect 9399 8676 9423 8678
rect 9479 8676 9503 8678
rect 9559 8676 9565 8678
rect 9257 8667 9565 8676
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8265 9444 8434
rect 9402 8256 9458 8265
rect 9402 8191 9458 8200
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9034 7984 9090 7993
rect 9034 7919 9090 7928
rect 9048 7886 9076 7919
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9048 7002 9076 7822
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9140 6866 9168 7686
rect 9257 7644 9565 7653
rect 9257 7642 9263 7644
rect 9319 7642 9343 7644
rect 9399 7642 9423 7644
rect 9479 7642 9503 7644
rect 9559 7642 9565 7644
rect 9319 7590 9321 7642
rect 9501 7590 9503 7642
rect 9257 7588 9263 7590
rect 9319 7588 9343 7590
rect 9399 7588 9423 7590
rect 9479 7588 9503 7590
rect 9559 7588 9565 7590
rect 9257 7579 9565 7588
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6866 9260 7142
rect 9416 6905 9444 7346
rect 9402 6896 9458 6905
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9220 6860 9272 6866
rect 9600 6866 9628 9318
rect 9402 6831 9458 6840
rect 9588 6860 9640 6866
rect 9220 6802 9272 6808
rect 9588 6802 9640 6808
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8484 6316 8536 6322
rect 8404 6276 8484 6304
rect 8404 5234 8432 6276
rect 8484 6258 8536 6264
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8220 4078 8248 4422
rect 8312 4185 8340 4626
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8024 4072 8076 4078
rect 8208 4072 8260 4078
rect 8076 4020 8156 4026
rect 8024 4014 8156 4020
rect 8208 4014 8260 4020
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3602 7604 3878
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7380 3528 7432 3534
rect 7208 3476 7380 3482
rect 7208 3470 7432 3476
rect 7208 3466 7420 3470
rect 7196 3460 7420 3466
rect 7248 3454 7420 3460
rect 7472 3460 7524 3466
rect 7196 3402 7248 3408
rect 7472 3402 7524 3408
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7072 3292 7380 3301
rect 7072 3290 7078 3292
rect 7134 3290 7158 3292
rect 7214 3290 7238 3292
rect 7294 3290 7318 3292
rect 7374 3290 7380 3292
rect 7134 3238 7136 3290
rect 7316 3238 7318 3290
rect 7072 3236 7078 3238
rect 7134 3236 7158 3238
rect 7214 3236 7238 3238
rect 7294 3236 7318 3238
rect 7374 3236 7380 3238
rect 7072 3227 7380 3236
rect 7484 3194 7512 3402
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7576 3074 7604 3402
rect 7484 3058 7604 3074
rect 7668 3058 7696 4014
rect 7944 3618 7972 4014
rect 8036 3998 8156 4014
rect 7944 3590 8064 3618
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7472 3052 7604 3058
rect 7524 3046 7604 3052
rect 7656 3052 7708 3058
rect 7472 2994 7524 3000
rect 7656 2994 7708 3000
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 6288 2446 6316 2790
rect 6412 2748 6720 2757
rect 6412 2746 6418 2748
rect 6474 2746 6498 2748
rect 6554 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6720 2748
rect 6474 2694 6476 2746
rect 6656 2694 6658 2746
rect 6412 2692 6418 2694
rect 6474 2692 6498 2694
rect 6554 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6720 2694
rect 6412 2683 6720 2692
rect 7760 2446 7788 3334
rect 7852 3194 7880 3470
rect 7944 3194 7972 3470
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8036 2990 8064 3590
rect 8128 3398 8156 3998
rect 8312 3534 8340 4014
rect 8404 3602 8432 5170
rect 8496 4622 8524 6122
rect 8597 6012 8905 6021
rect 8597 6010 8603 6012
rect 8659 6010 8683 6012
rect 8739 6010 8763 6012
rect 8819 6010 8843 6012
rect 8899 6010 8905 6012
rect 8659 5958 8661 6010
rect 8841 5958 8843 6010
rect 8597 5956 8603 5958
rect 8659 5956 8683 5958
rect 8739 5956 8763 5958
rect 8819 5956 8843 5958
rect 8899 5956 8905 5958
rect 8597 5947 8905 5956
rect 8956 5914 8984 6666
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5234 8984 5510
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8597 4924 8905 4933
rect 8597 4922 8603 4924
rect 8659 4922 8683 4924
rect 8739 4922 8763 4924
rect 8819 4922 8843 4924
rect 8899 4922 8905 4924
rect 8659 4870 8661 4922
rect 8841 4870 8843 4922
rect 8597 4868 8603 4870
rect 8659 4868 8683 4870
rect 8739 4868 8763 4870
rect 8819 4868 8843 4870
rect 8899 4868 8905 4870
rect 8597 4859 8905 4868
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8956 3942 8984 5170
rect 9140 4622 9168 6598
rect 9257 6556 9565 6565
rect 9257 6554 9263 6556
rect 9319 6554 9343 6556
rect 9399 6554 9423 6556
rect 9479 6554 9503 6556
rect 9559 6554 9565 6556
rect 9319 6502 9321 6554
rect 9501 6502 9503 6554
rect 9257 6500 9263 6502
rect 9319 6500 9343 6502
rect 9399 6500 9423 6502
rect 9479 6500 9503 6502
rect 9559 6500 9565 6502
rect 9257 6491 9565 6500
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5642 9260 6190
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9257 5468 9565 5477
rect 9257 5466 9263 5468
rect 9319 5466 9343 5468
rect 9399 5466 9423 5468
rect 9479 5466 9503 5468
rect 9559 5466 9565 5468
rect 9319 5414 9321 5466
rect 9501 5414 9503 5466
rect 9257 5412 9263 5414
rect 9319 5412 9343 5414
rect 9399 5412 9423 5414
rect 9479 5412 9503 5414
rect 9559 5412 9565 5414
rect 9257 5403 9565 5412
rect 9586 4856 9642 4865
rect 9586 4791 9642 4800
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9257 4380 9565 4389
rect 9257 4378 9263 4380
rect 9319 4378 9343 4380
rect 9399 4378 9423 4380
rect 9479 4378 9503 4380
rect 9559 4378 9565 4380
rect 9319 4326 9321 4378
rect 9501 4326 9503 4378
rect 9257 4324 9263 4326
rect 9319 4324 9343 4326
rect 9399 4324 9423 4326
rect 9479 4324 9503 4326
rect 9559 4324 9565 4326
rect 9257 4315 9565 4324
rect 9600 4146 9628 4791
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9692 4078 9720 4490
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8597 3836 8905 3845
rect 8597 3834 8603 3836
rect 8659 3834 8683 3836
rect 8739 3834 8763 3836
rect 8819 3834 8843 3836
rect 8899 3834 8905 3836
rect 8659 3782 8661 3834
rect 8841 3782 8843 3834
rect 8597 3780 8603 3782
rect 8659 3780 8683 3782
rect 8739 3780 8763 3782
rect 8819 3780 8843 3782
rect 8899 3780 8905 3782
rect 8597 3771 8905 3780
rect 9692 3602 9720 4014
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 9048 3126 9076 3402
rect 9257 3292 9565 3301
rect 9257 3290 9263 3292
rect 9319 3290 9343 3292
rect 9399 3290 9423 3292
rect 9479 3290 9503 3292
rect 9559 3290 9565 3292
rect 9319 3238 9321 3290
rect 9501 3238 9503 3290
rect 9257 3236 9263 3238
rect 9319 3236 9343 3238
rect 9399 3236 9423 3238
rect 9479 3236 9503 3238
rect 9559 3236 9565 3238
rect 9257 3227 9565 3236
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7852 2446 7880 2858
rect 8036 2650 8064 2926
rect 8312 2650 8340 2926
rect 8588 2854 8616 2994
rect 8576 2848 8628 2854
rect 8496 2808 8576 2836
rect 8496 2650 8524 2808
rect 8576 2790 8628 2796
rect 8597 2748 8905 2757
rect 8597 2746 8603 2748
rect 8659 2746 8683 2748
rect 8739 2746 8763 2748
rect 8819 2746 8843 2748
rect 8899 2746 8905 2748
rect 8659 2694 8661 2746
rect 8841 2694 8843 2746
rect 8597 2692 8603 2694
rect 8659 2692 8683 2694
rect 8739 2692 8763 2694
rect 8819 2692 8843 2694
rect 8899 2692 8905 2694
rect 8597 2683 8905 2692
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 2702 2204 3010 2213
rect 2702 2202 2708 2204
rect 2764 2202 2788 2204
rect 2844 2202 2868 2204
rect 2924 2202 2948 2204
rect 3004 2202 3010 2204
rect 2764 2150 2766 2202
rect 2946 2150 2948 2202
rect 2702 2148 2708 2150
rect 2764 2148 2788 2150
rect 2844 2148 2868 2150
rect 2924 2148 2948 2150
rect 3004 2148 3010 2150
rect 2702 2139 3010 2148
rect 3252 800 3280 2382
rect 3896 800 3924 2382
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4540 800 4568 2314
rect 4887 2204 5195 2213
rect 4887 2202 4893 2204
rect 4949 2202 4973 2204
rect 5029 2202 5053 2204
rect 5109 2202 5133 2204
rect 5189 2202 5195 2204
rect 4949 2150 4951 2202
rect 5131 2150 5133 2202
rect 4887 2148 4893 2150
rect 4949 2148 4973 2150
rect 5029 2148 5053 2150
rect 5109 2148 5133 2150
rect 5189 2148 5195 2150
rect 4887 2139 5195 2148
rect 5276 1306 5304 2382
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 5828 800 5856 2314
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 6932 1170 6960 2246
rect 7072 2204 7380 2213
rect 7072 2202 7078 2204
rect 7134 2202 7158 2204
rect 7214 2202 7238 2204
rect 7294 2202 7318 2204
rect 7374 2202 7380 2204
rect 7134 2150 7136 2202
rect 7316 2150 7318 2202
rect 7072 2148 7078 2150
rect 7134 2148 7158 2150
rect 7214 2148 7238 2150
rect 7294 2148 7318 2150
rect 7374 2148 7380 2150
rect 7072 2139 7380 2148
rect 6932 1142 7144 1170
rect 7116 800 7144 1142
rect 7760 800 7788 2246
rect 8404 800 8432 2382
rect 9257 2204 9565 2213
rect 9257 2202 9263 2204
rect 9319 2202 9343 2204
rect 9399 2202 9423 2204
rect 9479 2202 9503 2204
rect 9559 2202 9565 2204
rect 9319 2150 9321 2202
rect 9501 2150 9503 2202
rect 9257 2148 9263 2150
rect 9319 2148 9343 2150
rect 9399 2148 9423 2150
rect 9479 2148 9503 2150
rect 9559 2148 9565 2150
rect 9257 2139 9565 2148
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< via2 >>
rect 2708 10906 2764 10908
rect 2788 10906 2844 10908
rect 2868 10906 2924 10908
rect 2948 10906 3004 10908
rect 2708 10854 2754 10906
rect 2754 10854 2764 10906
rect 2788 10854 2818 10906
rect 2818 10854 2830 10906
rect 2830 10854 2844 10906
rect 2868 10854 2882 10906
rect 2882 10854 2894 10906
rect 2894 10854 2924 10906
rect 2948 10854 2958 10906
rect 2958 10854 3004 10906
rect 2708 10852 2764 10854
rect 2788 10852 2844 10854
rect 2868 10852 2924 10854
rect 2948 10852 3004 10854
rect 4893 10906 4949 10908
rect 4973 10906 5029 10908
rect 5053 10906 5109 10908
rect 5133 10906 5189 10908
rect 4893 10854 4939 10906
rect 4939 10854 4949 10906
rect 4973 10854 5003 10906
rect 5003 10854 5015 10906
rect 5015 10854 5029 10906
rect 5053 10854 5067 10906
rect 5067 10854 5079 10906
rect 5079 10854 5109 10906
rect 5133 10854 5143 10906
rect 5143 10854 5189 10906
rect 4893 10852 4949 10854
rect 4973 10852 5029 10854
rect 5053 10852 5109 10854
rect 5133 10852 5189 10854
rect 2048 10362 2104 10364
rect 2128 10362 2184 10364
rect 2208 10362 2264 10364
rect 2288 10362 2344 10364
rect 2048 10310 2094 10362
rect 2094 10310 2104 10362
rect 2128 10310 2158 10362
rect 2158 10310 2170 10362
rect 2170 10310 2184 10362
rect 2208 10310 2222 10362
rect 2222 10310 2234 10362
rect 2234 10310 2264 10362
rect 2288 10310 2298 10362
rect 2298 10310 2344 10362
rect 2048 10308 2104 10310
rect 2128 10308 2184 10310
rect 2208 10308 2264 10310
rect 2288 10308 2344 10310
rect 1398 9560 1454 9616
rect 2708 9818 2764 9820
rect 2788 9818 2844 9820
rect 2868 9818 2924 9820
rect 2948 9818 3004 9820
rect 2708 9766 2754 9818
rect 2754 9766 2764 9818
rect 2788 9766 2818 9818
rect 2818 9766 2830 9818
rect 2830 9766 2844 9818
rect 2868 9766 2882 9818
rect 2882 9766 2894 9818
rect 2894 9766 2924 9818
rect 2948 9766 2958 9818
rect 2958 9766 3004 9818
rect 2708 9764 2764 9766
rect 2788 9764 2844 9766
rect 2868 9764 2924 9766
rect 2948 9764 3004 9766
rect 7078 10906 7134 10908
rect 7158 10906 7214 10908
rect 7238 10906 7294 10908
rect 7318 10906 7374 10908
rect 7078 10854 7124 10906
rect 7124 10854 7134 10906
rect 7158 10854 7188 10906
rect 7188 10854 7200 10906
rect 7200 10854 7214 10906
rect 7238 10854 7252 10906
rect 7252 10854 7264 10906
rect 7264 10854 7294 10906
rect 7318 10854 7328 10906
rect 7328 10854 7374 10906
rect 7078 10852 7134 10854
rect 7158 10852 7214 10854
rect 7238 10852 7294 10854
rect 7318 10852 7374 10854
rect 4233 10362 4289 10364
rect 4313 10362 4369 10364
rect 4393 10362 4449 10364
rect 4473 10362 4529 10364
rect 4233 10310 4279 10362
rect 4279 10310 4289 10362
rect 4313 10310 4343 10362
rect 4343 10310 4355 10362
rect 4355 10310 4369 10362
rect 4393 10310 4407 10362
rect 4407 10310 4419 10362
rect 4419 10310 4449 10362
rect 4473 10310 4483 10362
rect 4483 10310 4529 10362
rect 4233 10308 4289 10310
rect 4313 10308 4369 10310
rect 4393 10308 4449 10310
rect 4473 10308 4529 10310
rect 2048 9274 2104 9276
rect 2128 9274 2184 9276
rect 2208 9274 2264 9276
rect 2288 9274 2344 9276
rect 2048 9222 2094 9274
rect 2094 9222 2104 9274
rect 2128 9222 2158 9274
rect 2158 9222 2170 9274
rect 2170 9222 2184 9274
rect 2208 9222 2222 9274
rect 2222 9222 2234 9274
rect 2234 9222 2264 9274
rect 2288 9222 2298 9274
rect 2298 9222 2344 9274
rect 2048 9220 2104 9222
rect 2128 9220 2184 9222
rect 2208 9220 2264 9222
rect 2288 9220 2344 9222
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 846 7656 902 7712
rect 4233 9274 4289 9276
rect 4313 9274 4369 9276
rect 4393 9274 4449 9276
rect 4473 9274 4529 9276
rect 4233 9222 4279 9274
rect 4279 9222 4289 9274
rect 4313 9222 4343 9274
rect 4343 9222 4355 9274
rect 4355 9222 4369 9274
rect 4393 9222 4407 9274
rect 4407 9222 4419 9274
rect 4419 9222 4449 9274
rect 4473 9222 4483 9274
rect 4483 9222 4529 9274
rect 4233 9220 4289 9222
rect 4313 9220 4369 9222
rect 4393 9220 4449 9222
rect 4473 9220 4529 9222
rect 4893 9818 4949 9820
rect 4973 9818 5029 9820
rect 5053 9818 5109 9820
rect 5133 9818 5189 9820
rect 4893 9766 4939 9818
rect 4939 9766 4949 9818
rect 4973 9766 5003 9818
rect 5003 9766 5015 9818
rect 5015 9766 5029 9818
rect 5053 9766 5067 9818
rect 5067 9766 5079 9818
rect 5079 9766 5109 9818
rect 5133 9766 5143 9818
rect 5143 9766 5189 9818
rect 4893 9764 4949 9766
rect 4973 9764 5029 9766
rect 5053 9764 5109 9766
rect 5133 9764 5189 9766
rect 2708 8730 2764 8732
rect 2788 8730 2844 8732
rect 2868 8730 2924 8732
rect 2948 8730 3004 8732
rect 2708 8678 2754 8730
rect 2754 8678 2764 8730
rect 2788 8678 2818 8730
rect 2818 8678 2830 8730
rect 2830 8678 2844 8730
rect 2868 8678 2882 8730
rect 2882 8678 2894 8730
rect 2894 8678 2924 8730
rect 2948 8678 2958 8730
rect 2958 8678 3004 8730
rect 2708 8676 2764 8678
rect 2788 8676 2844 8678
rect 2868 8676 2924 8678
rect 2948 8676 3004 8678
rect 2048 8186 2104 8188
rect 2128 8186 2184 8188
rect 2208 8186 2264 8188
rect 2288 8186 2344 8188
rect 2048 8134 2094 8186
rect 2094 8134 2104 8186
rect 2128 8134 2158 8186
rect 2158 8134 2170 8186
rect 2170 8134 2184 8186
rect 2208 8134 2222 8186
rect 2222 8134 2234 8186
rect 2234 8134 2264 8186
rect 2288 8134 2298 8186
rect 2298 8134 2344 8186
rect 2048 8132 2104 8134
rect 2128 8132 2184 8134
rect 2208 8132 2264 8134
rect 2288 8132 2344 8134
rect 1490 6840 1546 6896
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 1214 4820 1270 4856
rect 1214 4800 1216 4820
rect 1216 4800 1268 4820
rect 1268 4800 1270 4820
rect 2048 7098 2104 7100
rect 2128 7098 2184 7100
rect 2208 7098 2264 7100
rect 2288 7098 2344 7100
rect 2048 7046 2094 7098
rect 2094 7046 2104 7098
rect 2128 7046 2158 7098
rect 2158 7046 2170 7098
rect 2170 7046 2184 7098
rect 2208 7046 2222 7098
rect 2222 7046 2234 7098
rect 2234 7046 2264 7098
rect 2288 7046 2298 7098
rect 2298 7046 2344 7098
rect 2048 7044 2104 7046
rect 2128 7044 2184 7046
rect 2208 7044 2264 7046
rect 2288 7044 2344 7046
rect 2708 7642 2764 7644
rect 2788 7642 2844 7644
rect 2868 7642 2924 7644
rect 2948 7642 3004 7644
rect 2708 7590 2754 7642
rect 2754 7590 2764 7642
rect 2788 7590 2818 7642
rect 2818 7590 2830 7642
rect 2830 7590 2844 7642
rect 2868 7590 2882 7642
rect 2882 7590 2894 7642
rect 2894 7590 2924 7642
rect 2948 7590 2958 7642
rect 2958 7590 3004 7642
rect 2708 7588 2764 7590
rect 2788 7588 2844 7590
rect 2868 7588 2924 7590
rect 2948 7588 3004 7590
rect 4893 8730 4949 8732
rect 4973 8730 5029 8732
rect 5053 8730 5109 8732
rect 5133 8730 5189 8732
rect 4893 8678 4939 8730
rect 4939 8678 4949 8730
rect 4973 8678 5003 8730
rect 5003 8678 5015 8730
rect 5015 8678 5029 8730
rect 5053 8678 5067 8730
rect 5067 8678 5079 8730
rect 5079 8678 5109 8730
rect 5133 8678 5143 8730
rect 5143 8678 5189 8730
rect 4893 8676 4949 8678
rect 4973 8676 5029 8678
rect 5053 8676 5109 8678
rect 5133 8676 5189 8678
rect 4233 8186 4289 8188
rect 4313 8186 4369 8188
rect 4393 8186 4449 8188
rect 4473 8186 4529 8188
rect 4233 8134 4279 8186
rect 4279 8134 4289 8186
rect 4313 8134 4343 8186
rect 4343 8134 4355 8186
rect 4355 8134 4369 8186
rect 4393 8134 4407 8186
rect 4407 8134 4419 8186
rect 4419 8134 4449 8186
rect 4473 8134 4483 8186
rect 4483 8134 4529 8186
rect 4233 8132 4289 8134
rect 4313 8132 4369 8134
rect 4393 8132 4449 8134
rect 4473 8132 4529 8134
rect 4893 7642 4949 7644
rect 4973 7642 5029 7644
rect 5053 7642 5109 7644
rect 5133 7642 5189 7644
rect 4893 7590 4939 7642
rect 4939 7590 4949 7642
rect 4973 7590 5003 7642
rect 5003 7590 5015 7642
rect 5015 7590 5029 7642
rect 5053 7590 5067 7642
rect 5067 7590 5079 7642
rect 5079 7590 5109 7642
rect 5133 7590 5143 7642
rect 5143 7590 5189 7642
rect 4893 7588 4949 7590
rect 4973 7588 5029 7590
rect 5053 7588 5109 7590
rect 5133 7588 5189 7590
rect 4233 7098 4289 7100
rect 4313 7098 4369 7100
rect 4393 7098 4449 7100
rect 4473 7098 4529 7100
rect 4233 7046 4279 7098
rect 4279 7046 4289 7098
rect 4313 7046 4343 7098
rect 4343 7046 4355 7098
rect 4355 7046 4369 7098
rect 4393 7046 4407 7098
rect 4407 7046 4419 7098
rect 4419 7046 4449 7098
rect 4473 7046 4483 7098
rect 4483 7046 4529 7098
rect 4233 7044 4289 7046
rect 4313 7044 4369 7046
rect 4393 7044 4449 7046
rect 4473 7044 4529 7046
rect 1398 5480 1454 5536
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 2048 6010 2104 6012
rect 2128 6010 2184 6012
rect 2208 6010 2264 6012
rect 2288 6010 2344 6012
rect 2048 5958 2094 6010
rect 2094 5958 2104 6010
rect 2128 5958 2158 6010
rect 2158 5958 2170 6010
rect 2170 5958 2184 6010
rect 2208 5958 2222 6010
rect 2222 5958 2234 6010
rect 2234 5958 2264 6010
rect 2288 5958 2298 6010
rect 2298 5958 2344 6010
rect 2048 5956 2104 5958
rect 2128 5956 2184 5958
rect 2208 5956 2264 5958
rect 2288 5956 2344 5958
rect 2048 4922 2104 4924
rect 2128 4922 2184 4924
rect 2208 4922 2264 4924
rect 2288 4922 2344 4924
rect 2048 4870 2094 4922
rect 2094 4870 2104 4922
rect 2128 4870 2158 4922
rect 2158 4870 2170 4922
rect 2170 4870 2184 4922
rect 2208 4870 2222 4922
rect 2222 4870 2234 4922
rect 2234 4870 2264 4922
rect 2288 4870 2298 4922
rect 2298 4870 2344 4922
rect 2048 4868 2104 4870
rect 2128 4868 2184 4870
rect 2208 4868 2264 4870
rect 2288 4868 2344 4870
rect 2708 6554 2764 6556
rect 2788 6554 2844 6556
rect 2868 6554 2924 6556
rect 2948 6554 3004 6556
rect 2708 6502 2754 6554
rect 2754 6502 2764 6554
rect 2788 6502 2818 6554
rect 2818 6502 2830 6554
rect 2830 6502 2844 6554
rect 2868 6502 2882 6554
rect 2882 6502 2894 6554
rect 2894 6502 2924 6554
rect 2948 6502 2958 6554
rect 2958 6502 3004 6554
rect 2708 6500 2764 6502
rect 2788 6500 2844 6502
rect 2868 6500 2924 6502
rect 2948 6500 3004 6502
rect 2708 5466 2764 5468
rect 2788 5466 2844 5468
rect 2868 5466 2924 5468
rect 2948 5466 3004 5468
rect 2708 5414 2754 5466
rect 2754 5414 2764 5466
rect 2788 5414 2818 5466
rect 2818 5414 2830 5466
rect 2830 5414 2844 5466
rect 2868 5414 2882 5466
rect 2882 5414 2894 5466
rect 2894 5414 2924 5466
rect 2948 5414 2958 5466
rect 2958 5414 3004 5466
rect 2708 5412 2764 5414
rect 2788 5412 2844 5414
rect 2868 5412 2924 5414
rect 2948 5412 3004 5414
rect 4233 6010 4289 6012
rect 4313 6010 4369 6012
rect 4393 6010 4449 6012
rect 4473 6010 4529 6012
rect 4233 5958 4279 6010
rect 4279 5958 4289 6010
rect 4313 5958 4343 6010
rect 4343 5958 4355 6010
rect 4355 5958 4369 6010
rect 4393 5958 4407 6010
rect 4407 5958 4419 6010
rect 4419 5958 4449 6010
rect 4473 5958 4483 6010
rect 4483 5958 4529 6010
rect 4233 5956 4289 5958
rect 4313 5956 4369 5958
rect 4393 5956 4449 5958
rect 4473 5956 4529 5958
rect 2594 5244 2596 5264
rect 2596 5244 2648 5264
rect 2648 5244 2650 5264
rect 2594 5208 2650 5244
rect 2708 4378 2764 4380
rect 2788 4378 2844 4380
rect 2868 4378 2924 4380
rect 2948 4378 3004 4380
rect 2708 4326 2754 4378
rect 2754 4326 2764 4378
rect 2788 4326 2818 4378
rect 2818 4326 2830 4378
rect 2830 4326 2844 4378
rect 2868 4326 2882 4378
rect 2882 4326 2894 4378
rect 2894 4326 2924 4378
rect 2948 4326 2958 4378
rect 2958 4326 3004 4378
rect 2708 4324 2764 4326
rect 2788 4324 2844 4326
rect 2868 4324 2924 4326
rect 2948 4324 3004 4326
rect 2048 3834 2104 3836
rect 2128 3834 2184 3836
rect 2208 3834 2264 3836
rect 2288 3834 2344 3836
rect 2048 3782 2094 3834
rect 2094 3782 2104 3834
rect 2128 3782 2158 3834
rect 2158 3782 2170 3834
rect 2170 3782 2184 3834
rect 2208 3782 2222 3834
rect 2222 3782 2234 3834
rect 2234 3782 2264 3834
rect 2288 3782 2298 3834
rect 2298 3782 2344 3834
rect 2048 3780 2104 3782
rect 2128 3780 2184 3782
rect 2208 3780 2264 3782
rect 2288 3780 2344 3782
rect 2708 3290 2764 3292
rect 2788 3290 2844 3292
rect 2868 3290 2924 3292
rect 2948 3290 3004 3292
rect 2708 3238 2754 3290
rect 2754 3238 2764 3290
rect 2788 3238 2818 3290
rect 2818 3238 2830 3290
rect 2830 3238 2844 3290
rect 2868 3238 2882 3290
rect 2882 3238 2894 3290
rect 2894 3238 2924 3290
rect 2948 3238 2958 3290
rect 2958 3238 3004 3290
rect 2708 3236 2764 3238
rect 2788 3236 2844 3238
rect 2868 3236 2924 3238
rect 2948 3236 3004 3238
rect 2048 2746 2104 2748
rect 2128 2746 2184 2748
rect 2208 2746 2264 2748
rect 2288 2746 2344 2748
rect 2048 2694 2094 2746
rect 2094 2694 2104 2746
rect 2128 2694 2158 2746
rect 2158 2694 2170 2746
rect 2170 2694 2184 2746
rect 2208 2694 2222 2746
rect 2222 2694 2234 2746
rect 2234 2694 2264 2746
rect 2288 2694 2298 2746
rect 2298 2694 2344 2746
rect 2048 2692 2104 2694
rect 2128 2692 2184 2694
rect 2208 2692 2264 2694
rect 2288 2692 2344 2694
rect 4526 5092 4582 5128
rect 4526 5072 4528 5092
rect 4528 5072 4580 5092
rect 4580 5072 4582 5092
rect 4233 4922 4289 4924
rect 4313 4922 4369 4924
rect 4393 4922 4449 4924
rect 4473 4922 4529 4924
rect 4233 4870 4279 4922
rect 4279 4870 4289 4922
rect 4313 4870 4343 4922
rect 4343 4870 4355 4922
rect 4355 4870 4369 4922
rect 4393 4870 4407 4922
rect 4407 4870 4419 4922
rect 4419 4870 4449 4922
rect 4473 4870 4483 4922
rect 4483 4870 4529 4922
rect 4233 4868 4289 4870
rect 4313 4868 4369 4870
rect 4393 4868 4449 4870
rect 4473 4868 4529 4870
rect 6418 10362 6474 10364
rect 6498 10362 6554 10364
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6418 10310 6464 10362
rect 6464 10310 6474 10362
rect 6498 10310 6528 10362
rect 6528 10310 6540 10362
rect 6540 10310 6554 10362
rect 6578 10310 6592 10362
rect 6592 10310 6604 10362
rect 6604 10310 6634 10362
rect 6658 10310 6668 10362
rect 6668 10310 6714 10362
rect 6418 10308 6474 10310
rect 6498 10308 6554 10310
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 7078 9818 7134 9820
rect 7158 9818 7214 9820
rect 7238 9818 7294 9820
rect 7318 9818 7374 9820
rect 7078 9766 7124 9818
rect 7124 9766 7134 9818
rect 7158 9766 7188 9818
rect 7188 9766 7200 9818
rect 7200 9766 7214 9818
rect 7238 9766 7252 9818
rect 7252 9766 7264 9818
rect 7264 9766 7294 9818
rect 7318 9766 7328 9818
rect 7328 9766 7374 9818
rect 7078 9764 7134 9766
rect 7158 9764 7214 9766
rect 7238 9764 7294 9766
rect 7318 9764 7374 9766
rect 6418 9274 6474 9276
rect 6498 9274 6554 9276
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6418 9222 6464 9274
rect 6464 9222 6474 9274
rect 6498 9222 6528 9274
rect 6528 9222 6540 9274
rect 6540 9222 6554 9274
rect 6578 9222 6592 9274
rect 6592 9222 6604 9274
rect 6604 9222 6634 9274
rect 6658 9222 6668 9274
rect 6668 9222 6714 9274
rect 6418 9220 6474 9222
rect 6498 9220 6554 9222
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 7078 8730 7134 8732
rect 7158 8730 7214 8732
rect 7238 8730 7294 8732
rect 7318 8730 7374 8732
rect 7078 8678 7124 8730
rect 7124 8678 7134 8730
rect 7158 8678 7188 8730
rect 7188 8678 7200 8730
rect 7200 8678 7214 8730
rect 7238 8678 7252 8730
rect 7252 8678 7264 8730
rect 7264 8678 7294 8730
rect 7318 8678 7328 8730
rect 7328 8678 7374 8730
rect 7078 8676 7134 8678
rect 7158 8676 7214 8678
rect 7238 8676 7294 8678
rect 7318 8676 7374 8678
rect 4893 6554 4949 6556
rect 4973 6554 5029 6556
rect 5053 6554 5109 6556
rect 5133 6554 5189 6556
rect 4893 6502 4939 6554
rect 4939 6502 4949 6554
rect 4973 6502 5003 6554
rect 5003 6502 5015 6554
rect 5015 6502 5029 6554
rect 5053 6502 5067 6554
rect 5067 6502 5079 6554
rect 5079 6502 5109 6554
rect 5133 6502 5143 6554
rect 5143 6502 5189 6554
rect 4893 6500 4949 6502
rect 4973 6500 5029 6502
rect 5053 6500 5109 6502
rect 5133 6500 5189 6502
rect 6418 8186 6474 8188
rect 6498 8186 6554 8188
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6418 8134 6464 8186
rect 6464 8134 6474 8186
rect 6498 8134 6528 8186
rect 6528 8134 6540 8186
rect 6540 8134 6554 8186
rect 6578 8134 6592 8186
rect 6592 8134 6604 8186
rect 6604 8134 6634 8186
rect 6658 8134 6668 8186
rect 6668 8134 6714 8186
rect 6418 8132 6474 8134
rect 6498 8132 6554 8134
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 7102 8472 7158 8528
rect 7378 7928 7434 7984
rect 6418 7098 6474 7100
rect 6498 7098 6554 7100
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6418 7046 6464 7098
rect 6464 7046 6474 7098
rect 6498 7046 6528 7098
rect 6528 7046 6540 7098
rect 6540 7046 6554 7098
rect 6578 7046 6592 7098
rect 6592 7046 6604 7098
rect 6604 7046 6634 7098
rect 6658 7046 6668 7098
rect 6668 7046 6714 7098
rect 6418 7044 6474 7046
rect 6498 7044 6554 7046
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 7078 7642 7134 7644
rect 7158 7642 7214 7644
rect 7238 7642 7294 7644
rect 7318 7642 7374 7644
rect 7078 7590 7124 7642
rect 7124 7590 7134 7642
rect 7158 7590 7188 7642
rect 7188 7590 7200 7642
rect 7200 7590 7214 7642
rect 7238 7590 7252 7642
rect 7252 7590 7264 7642
rect 7264 7590 7294 7642
rect 7318 7590 7328 7642
rect 7328 7590 7374 7642
rect 7078 7588 7134 7590
rect 7158 7588 7214 7590
rect 7238 7588 7294 7590
rect 7318 7588 7374 7590
rect 7378 7384 7434 7440
rect 7654 7928 7710 7984
rect 4893 5466 4949 5468
rect 4973 5466 5029 5468
rect 5053 5466 5109 5468
rect 5133 5466 5189 5468
rect 4893 5414 4939 5466
rect 4939 5414 4949 5466
rect 4973 5414 5003 5466
rect 5003 5414 5015 5466
rect 5015 5414 5029 5466
rect 5053 5414 5067 5466
rect 5067 5414 5079 5466
rect 5079 5414 5109 5466
rect 5133 5414 5143 5466
rect 5143 5414 5189 5466
rect 4893 5412 4949 5414
rect 4973 5412 5029 5414
rect 5053 5412 5109 5414
rect 5133 5412 5189 5414
rect 5262 5244 5264 5264
rect 5264 5244 5316 5264
rect 5316 5244 5318 5264
rect 5262 5208 5318 5244
rect 4710 5072 4766 5128
rect 4233 3834 4289 3836
rect 4313 3834 4369 3836
rect 4393 3834 4449 3836
rect 4473 3834 4529 3836
rect 4233 3782 4279 3834
rect 4279 3782 4289 3834
rect 4313 3782 4343 3834
rect 4343 3782 4355 3834
rect 4355 3782 4369 3834
rect 4393 3782 4407 3834
rect 4407 3782 4419 3834
rect 4419 3782 4449 3834
rect 4473 3782 4483 3834
rect 4483 3782 4529 3834
rect 4233 3780 4289 3782
rect 4313 3780 4369 3782
rect 4393 3780 4449 3782
rect 4473 3780 4529 3782
rect 4233 2746 4289 2748
rect 4313 2746 4369 2748
rect 4393 2746 4449 2748
rect 4473 2746 4529 2748
rect 4233 2694 4279 2746
rect 4279 2694 4289 2746
rect 4313 2694 4343 2746
rect 4343 2694 4355 2746
rect 4355 2694 4369 2746
rect 4393 2694 4407 2746
rect 4407 2694 4419 2746
rect 4419 2694 4449 2746
rect 4473 2694 4483 2746
rect 4483 2694 4529 2746
rect 4233 2692 4289 2694
rect 4313 2692 4369 2694
rect 4393 2692 4449 2694
rect 4473 2692 4529 2694
rect 4893 4378 4949 4380
rect 4973 4378 5029 4380
rect 5053 4378 5109 4380
rect 5133 4378 5189 4380
rect 4893 4326 4939 4378
rect 4939 4326 4949 4378
rect 4973 4326 5003 4378
rect 5003 4326 5015 4378
rect 5015 4326 5029 4378
rect 5053 4326 5067 4378
rect 5067 4326 5079 4378
rect 5079 4326 5109 4378
rect 5133 4326 5143 4378
rect 5143 4326 5189 4378
rect 4893 4324 4949 4326
rect 4973 4324 5029 4326
rect 5053 4324 5109 4326
rect 5133 4324 5189 4326
rect 4893 3290 4949 3292
rect 4973 3290 5029 3292
rect 5053 3290 5109 3292
rect 5133 3290 5189 3292
rect 4893 3238 4939 3290
rect 4939 3238 4949 3290
rect 4973 3238 5003 3290
rect 5003 3238 5015 3290
rect 5015 3238 5029 3290
rect 5053 3238 5067 3290
rect 5067 3238 5079 3290
rect 5079 3238 5109 3290
rect 5133 3238 5143 3290
rect 5143 3238 5189 3290
rect 4893 3236 4949 3238
rect 4973 3236 5029 3238
rect 5053 3236 5109 3238
rect 5133 3236 5189 3238
rect 7078 6554 7134 6556
rect 7158 6554 7214 6556
rect 7238 6554 7294 6556
rect 7318 6554 7374 6556
rect 7078 6502 7124 6554
rect 7124 6502 7134 6554
rect 7158 6502 7188 6554
rect 7188 6502 7200 6554
rect 7200 6502 7214 6554
rect 7238 6502 7252 6554
rect 7252 6502 7264 6554
rect 7264 6502 7294 6554
rect 7318 6502 7328 6554
rect 7328 6502 7374 6554
rect 7078 6500 7134 6502
rect 7158 6500 7214 6502
rect 7238 6500 7294 6502
rect 7318 6500 7374 6502
rect 7470 6180 7526 6216
rect 7470 6160 7472 6180
rect 7472 6160 7524 6180
rect 7524 6160 7526 6180
rect 6418 6010 6474 6012
rect 6498 6010 6554 6012
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6418 5958 6464 6010
rect 6464 5958 6474 6010
rect 6498 5958 6528 6010
rect 6528 5958 6540 6010
rect 6540 5958 6554 6010
rect 6578 5958 6592 6010
rect 6592 5958 6604 6010
rect 6604 5958 6634 6010
rect 6658 5958 6668 6010
rect 6668 5958 6714 6010
rect 6418 5956 6474 5958
rect 6498 5956 6554 5958
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 9263 10906 9319 10908
rect 9343 10906 9399 10908
rect 9423 10906 9479 10908
rect 9503 10906 9559 10908
rect 9263 10854 9309 10906
rect 9309 10854 9319 10906
rect 9343 10854 9373 10906
rect 9373 10854 9385 10906
rect 9385 10854 9399 10906
rect 9423 10854 9437 10906
rect 9437 10854 9449 10906
rect 9449 10854 9479 10906
rect 9503 10854 9513 10906
rect 9513 10854 9559 10906
rect 9263 10852 9319 10854
rect 9343 10852 9399 10854
rect 9423 10852 9479 10854
rect 9503 10852 9559 10854
rect 8603 10362 8659 10364
rect 8683 10362 8739 10364
rect 8763 10362 8819 10364
rect 8843 10362 8899 10364
rect 8603 10310 8649 10362
rect 8649 10310 8659 10362
rect 8683 10310 8713 10362
rect 8713 10310 8725 10362
rect 8725 10310 8739 10362
rect 8763 10310 8777 10362
rect 8777 10310 8789 10362
rect 8789 10310 8819 10362
rect 8843 10310 8853 10362
rect 8853 10310 8899 10362
rect 8603 10308 8659 10310
rect 8683 10308 8739 10310
rect 8763 10308 8819 10310
rect 8843 10308 8899 10310
rect 8022 9444 8078 9480
rect 9263 9818 9319 9820
rect 9343 9818 9399 9820
rect 9423 9818 9479 9820
rect 9503 9818 9559 9820
rect 9263 9766 9309 9818
rect 9309 9766 9319 9818
rect 9343 9766 9373 9818
rect 9373 9766 9385 9818
rect 9385 9766 9399 9818
rect 9423 9766 9437 9818
rect 9437 9766 9449 9818
rect 9449 9766 9479 9818
rect 9503 9766 9513 9818
rect 9513 9766 9559 9818
rect 9263 9764 9319 9766
rect 9343 9764 9399 9766
rect 9423 9764 9479 9766
rect 9503 9764 9559 9766
rect 8022 9424 8024 9444
rect 8024 9424 8076 9444
rect 8076 9424 8078 9444
rect 8758 9460 8760 9480
rect 8760 9460 8812 9480
rect 8812 9460 8814 9480
rect 8758 9424 8814 9460
rect 8603 9274 8659 9276
rect 8683 9274 8739 9276
rect 8763 9274 8819 9276
rect 8843 9274 8899 9276
rect 8603 9222 8649 9274
rect 8649 9222 8659 9274
rect 8683 9222 8713 9274
rect 8713 9222 8725 9274
rect 8725 9222 8739 9274
rect 8763 9222 8777 9274
rect 8777 9222 8789 9274
rect 8789 9222 8819 9274
rect 8843 9222 8853 9274
rect 8853 9222 8899 9274
rect 8603 9220 8659 9222
rect 8683 9220 8739 9222
rect 8763 9220 8819 9222
rect 8843 9220 8899 9222
rect 8574 8472 8630 8528
rect 8603 8186 8659 8188
rect 8683 8186 8739 8188
rect 8763 8186 8819 8188
rect 8843 8186 8899 8188
rect 8603 8134 8649 8186
rect 8649 8134 8659 8186
rect 8683 8134 8713 8186
rect 8713 8134 8725 8186
rect 8725 8134 8739 8186
rect 8763 8134 8777 8186
rect 8777 8134 8789 8186
rect 8789 8134 8819 8186
rect 8843 8134 8853 8186
rect 8853 8134 8899 8186
rect 8603 8132 8659 8134
rect 8683 8132 8739 8134
rect 8763 8132 8819 8134
rect 8843 8132 8899 8134
rect 7078 5466 7134 5468
rect 7158 5466 7214 5468
rect 7238 5466 7294 5468
rect 7318 5466 7374 5468
rect 7078 5414 7124 5466
rect 7124 5414 7134 5466
rect 7158 5414 7188 5466
rect 7188 5414 7200 5466
rect 7200 5414 7214 5466
rect 7238 5414 7252 5466
rect 7252 5414 7264 5466
rect 7264 5414 7294 5466
rect 7318 5414 7328 5466
rect 7328 5414 7374 5466
rect 7078 5412 7134 5414
rect 7158 5412 7214 5414
rect 7238 5412 7294 5414
rect 7318 5412 7374 5414
rect 7194 5228 7250 5264
rect 7194 5208 7196 5228
rect 7196 5208 7248 5228
rect 7248 5208 7250 5228
rect 6418 4922 6474 4924
rect 6498 4922 6554 4924
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6418 4870 6464 4922
rect 6464 4870 6474 4922
rect 6498 4870 6528 4922
rect 6528 4870 6540 4922
rect 6540 4870 6554 4922
rect 6578 4870 6592 4922
rect 6592 4870 6604 4922
rect 6604 4870 6634 4922
rect 6658 4870 6668 4922
rect 6668 4870 6714 4922
rect 6418 4868 6474 4870
rect 6498 4868 6554 4870
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6418 3834 6474 3836
rect 6498 3834 6554 3836
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6418 3782 6464 3834
rect 6464 3782 6474 3834
rect 6498 3782 6528 3834
rect 6528 3782 6540 3834
rect 6540 3782 6554 3834
rect 6578 3782 6592 3834
rect 6592 3782 6604 3834
rect 6604 3782 6634 3834
rect 6658 3782 6668 3834
rect 6668 3782 6714 3834
rect 6418 3780 6474 3782
rect 6498 3780 6554 3782
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 7078 4378 7134 4380
rect 7158 4378 7214 4380
rect 7238 4378 7294 4380
rect 7318 4378 7374 4380
rect 7078 4326 7124 4378
rect 7124 4326 7134 4378
rect 7158 4326 7188 4378
rect 7188 4326 7200 4378
rect 7200 4326 7214 4378
rect 7238 4326 7252 4378
rect 7252 4326 7264 4378
rect 7264 4326 7294 4378
rect 7318 4326 7328 4378
rect 7328 4326 7374 4378
rect 7078 4324 7134 4326
rect 7158 4324 7214 4326
rect 7238 4324 7294 4326
rect 7318 4324 7374 4326
rect 8603 7098 8659 7100
rect 8683 7098 8739 7100
rect 8763 7098 8819 7100
rect 8843 7098 8899 7100
rect 8603 7046 8649 7098
rect 8649 7046 8659 7098
rect 8683 7046 8713 7098
rect 8713 7046 8725 7098
rect 8725 7046 8739 7098
rect 8763 7046 8777 7098
rect 8777 7046 8789 7098
rect 8789 7046 8819 7098
rect 8843 7046 8853 7098
rect 8853 7046 8899 7098
rect 8603 7044 8659 7046
rect 8683 7044 8739 7046
rect 8763 7044 8819 7046
rect 8843 7044 8899 7046
rect 9263 8730 9319 8732
rect 9343 8730 9399 8732
rect 9423 8730 9479 8732
rect 9503 8730 9559 8732
rect 9263 8678 9309 8730
rect 9309 8678 9319 8730
rect 9343 8678 9373 8730
rect 9373 8678 9385 8730
rect 9385 8678 9399 8730
rect 9423 8678 9437 8730
rect 9437 8678 9449 8730
rect 9449 8678 9479 8730
rect 9503 8678 9513 8730
rect 9513 8678 9559 8730
rect 9263 8676 9319 8678
rect 9343 8676 9399 8678
rect 9423 8676 9479 8678
rect 9503 8676 9559 8678
rect 9402 8200 9458 8256
rect 9034 7928 9090 7984
rect 9263 7642 9319 7644
rect 9343 7642 9399 7644
rect 9423 7642 9479 7644
rect 9503 7642 9559 7644
rect 9263 7590 9309 7642
rect 9309 7590 9319 7642
rect 9343 7590 9373 7642
rect 9373 7590 9385 7642
rect 9385 7590 9399 7642
rect 9423 7590 9437 7642
rect 9437 7590 9449 7642
rect 9449 7590 9479 7642
rect 9503 7590 9513 7642
rect 9513 7590 9559 7642
rect 9263 7588 9319 7590
rect 9343 7588 9399 7590
rect 9423 7588 9479 7590
rect 9503 7588 9559 7590
rect 9402 6840 9458 6896
rect 8298 4120 8354 4176
rect 7078 3290 7134 3292
rect 7158 3290 7214 3292
rect 7238 3290 7294 3292
rect 7318 3290 7374 3292
rect 7078 3238 7124 3290
rect 7124 3238 7134 3290
rect 7158 3238 7188 3290
rect 7188 3238 7200 3290
rect 7200 3238 7214 3290
rect 7238 3238 7252 3290
rect 7252 3238 7264 3290
rect 7264 3238 7294 3290
rect 7318 3238 7328 3290
rect 7328 3238 7374 3290
rect 7078 3236 7134 3238
rect 7158 3236 7214 3238
rect 7238 3236 7294 3238
rect 7318 3236 7374 3238
rect 6418 2746 6474 2748
rect 6498 2746 6554 2748
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6418 2694 6464 2746
rect 6464 2694 6474 2746
rect 6498 2694 6528 2746
rect 6528 2694 6540 2746
rect 6540 2694 6554 2746
rect 6578 2694 6592 2746
rect 6592 2694 6604 2746
rect 6604 2694 6634 2746
rect 6658 2694 6668 2746
rect 6668 2694 6714 2746
rect 6418 2692 6474 2694
rect 6498 2692 6554 2694
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 8603 6010 8659 6012
rect 8683 6010 8739 6012
rect 8763 6010 8819 6012
rect 8843 6010 8899 6012
rect 8603 5958 8649 6010
rect 8649 5958 8659 6010
rect 8683 5958 8713 6010
rect 8713 5958 8725 6010
rect 8725 5958 8739 6010
rect 8763 5958 8777 6010
rect 8777 5958 8789 6010
rect 8789 5958 8819 6010
rect 8843 5958 8853 6010
rect 8853 5958 8899 6010
rect 8603 5956 8659 5958
rect 8683 5956 8739 5958
rect 8763 5956 8819 5958
rect 8843 5956 8899 5958
rect 8603 4922 8659 4924
rect 8683 4922 8739 4924
rect 8763 4922 8819 4924
rect 8843 4922 8899 4924
rect 8603 4870 8649 4922
rect 8649 4870 8659 4922
rect 8683 4870 8713 4922
rect 8713 4870 8725 4922
rect 8725 4870 8739 4922
rect 8763 4870 8777 4922
rect 8777 4870 8789 4922
rect 8789 4870 8819 4922
rect 8843 4870 8853 4922
rect 8853 4870 8899 4922
rect 8603 4868 8659 4870
rect 8683 4868 8739 4870
rect 8763 4868 8819 4870
rect 8843 4868 8899 4870
rect 9263 6554 9319 6556
rect 9343 6554 9399 6556
rect 9423 6554 9479 6556
rect 9503 6554 9559 6556
rect 9263 6502 9309 6554
rect 9309 6502 9319 6554
rect 9343 6502 9373 6554
rect 9373 6502 9385 6554
rect 9385 6502 9399 6554
rect 9423 6502 9437 6554
rect 9437 6502 9449 6554
rect 9449 6502 9479 6554
rect 9503 6502 9513 6554
rect 9513 6502 9559 6554
rect 9263 6500 9319 6502
rect 9343 6500 9399 6502
rect 9423 6500 9479 6502
rect 9503 6500 9559 6502
rect 9263 5466 9319 5468
rect 9343 5466 9399 5468
rect 9423 5466 9479 5468
rect 9503 5466 9559 5468
rect 9263 5414 9309 5466
rect 9309 5414 9319 5466
rect 9343 5414 9373 5466
rect 9373 5414 9385 5466
rect 9385 5414 9399 5466
rect 9423 5414 9437 5466
rect 9437 5414 9449 5466
rect 9449 5414 9479 5466
rect 9503 5414 9513 5466
rect 9513 5414 9559 5466
rect 9263 5412 9319 5414
rect 9343 5412 9399 5414
rect 9423 5412 9479 5414
rect 9503 5412 9559 5414
rect 9586 4800 9642 4856
rect 9263 4378 9319 4380
rect 9343 4378 9399 4380
rect 9423 4378 9479 4380
rect 9503 4378 9559 4380
rect 9263 4326 9309 4378
rect 9309 4326 9319 4378
rect 9343 4326 9373 4378
rect 9373 4326 9385 4378
rect 9385 4326 9399 4378
rect 9423 4326 9437 4378
rect 9437 4326 9449 4378
rect 9449 4326 9479 4378
rect 9503 4326 9513 4378
rect 9513 4326 9559 4378
rect 9263 4324 9319 4326
rect 9343 4324 9399 4326
rect 9423 4324 9479 4326
rect 9503 4324 9559 4326
rect 8603 3834 8659 3836
rect 8683 3834 8739 3836
rect 8763 3834 8819 3836
rect 8843 3834 8899 3836
rect 8603 3782 8649 3834
rect 8649 3782 8659 3834
rect 8683 3782 8713 3834
rect 8713 3782 8725 3834
rect 8725 3782 8739 3834
rect 8763 3782 8777 3834
rect 8777 3782 8789 3834
rect 8789 3782 8819 3834
rect 8843 3782 8853 3834
rect 8853 3782 8899 3834
rect 8603 3780 8659 3782
rect 8683 3780 8739 3782
rect 8763 3780 8819 3782
rect 8843 3780 8899 3782
rect 9263 3290 9319 3292
rect 9343 3290 9399 3292
rect 9423 3290 9479 3292
rect 9503 3290 9559 3292
rect 9263 3238 9309 3290
rect 9309 3238 9319 3290
rect 9343 3238 9373 3290
rect 9373 3238 9385 3290
rect 9385 3238 9399 3290
rect 9423 3238 9437 3290
rect 9437 3238 9449 3290
rect 9449 3238 9479 3290
rect 9503 3238 9513 3290
rect 9513 3238 9559 3290
rect 9263 3236 9319 3238
rect 9343 3236 9399 3238
rect 9423 3236 9479 3238
rect 9503 3236 9559 3238
rect 8603 2746 8659 2748
rect 8683 2746 8739 2748
rect 8763 2746 8819 2748
rect 8843 2746 8899 2748
rect 8603 2694 8649 2746
rect 8649 2694 8659 2746
rect 8683 2694 8713 2746
rect 8713 2694 8725 2746
rect 8725 2694 8739 2746
rect 8763 2694 8777 2746
rect 8777 2694 8789 2746
rect 8789 2694 8819 2746
rect 8843 2694 8853 2746
rect 8853 2694 8899 2746
rect 8603 2692 8659 2694
rect 8683 2692 8739 2694
rect 8763 2692 8819 2694
rect 8843 2692 8899 2694
rect 2708 2202 2764 2204
rect 2788 2202 2844 2204
rect 2868 2202 2924 2204
rect 2948 2202 3004 2204
rect 2708 2150 2754 2202
rect 2754 2150 2764 2202
rect 2788 2150 2818 2202
rect 2818 2150 2830 2202
rect 2830 2150 2844 2202
rect 2868 2150 2882 2202
rect 2882 2150 2894 2202
rect 2894 2150 2924 2202
rect 2948 2150 2958 2202
rect 2958 2150 3004 2202
rect 2708 2148 2764 2150
rect 2788 2148 2844 2150
rect 2868 2148 2924 2150
rect 2948 2148 3004 2150
rect 4893 2202 4949 2204
rect 4973 2202 5029 2204
rect 5053 2202 5109 2204
rect 5133 2202 5189 2204
rect 4893 2150 4939 2202
rect 4939 2150 4949 2202
rect 4973 2150 5003 2202
rect 5003 2150 5015 2202
rect 5015 2150 5029 2202
rect 5053 2150 5067 2202
rect 5067 2150 5079 2202
rect 5079 2150 5109 2202
rect 5133 2150 5143 2202
rect 5143 2150 5189 2202
rect 4893 2148 4949 2150
rect 4973 2148 5029 2150
rect 5053 2148 5109 2150
rect 5133 2148 5189 2150
rect 7078 2202 7134 2204
rect 7158 2202 7214 2204
rect 7238 2202 7294 2204
rect 7318 2202 7374 2204
rect 7078 2150 7124 2202
rect 7124 2150 7134 2202
rect 7158 2150 7188 2202
rect 7188 2150 7200 2202
rect 7200 2150 7214 2202
rect 7238 2150 7252 2202
rect 7252 2150 7264 2202
rect 7264 2150 7294 2202
rect 7318 2150 7328 2202
rect 7328 2150 7374 2202
rect 7078 2148 7134 2150
rect 7158 2148 7214 2150
rect 7238 2148 7294 2150
rect 7318 2148 7374 2150
rect 9263 2202 9319 2204
rect 9343 2202 9399 2204
rect 9423 2202 9479 2204
rect 9503 2202 9559 2204
rect 9263 2150 9309 2202
rect 9309 2150 9319 2202
rect 9343 2150 9373 2202
rect 9373 2150 9385 2202
rect 9385 2150 9399 2202
rect 9423 2150 9437 2202
rect 9437 2150 9449 2202
rect 9449 2150 9479 2202
rect 9503 2150 9513 2202
rect 9513 2150 9559 2202
rect 9263 2148 9319 2150
rect 9343 2148 9399 2150
rect 9423 2148 9479 2150
rect 9503 2148 9559 2150
<< metal3 >>
rect 2698 10912 3014 10913
rect 2698 10848 2704 10912
rect 2768 10848 2784 10912
rect 2848 10848 2864 10912
rect 2928 10848 2944 10912
rect 3008 10848 3014 10912
rect 2698 10847 3014 10848
rect 4883 10912 5199 10913
rect 4883 10848 4889 10912
rect 4953 10848 4969 10912
rect 5033 10848 5049 10912
rect 5113 10848 5129 10912
rect 5193 10848 5199 10912
rect 4883 10847 5199 10848
rect 7068 10912 7384 10913
rect 7068 10848 7074 10912
rect 7138 10848 7154 10912
rect 7218 10848 7234 10912
rect 7298 10848 7314 10912
rect 7378 10848 7384 10912
rect 7068 10847 7384 10848
rect 9253 10912 9569 10913
rect 9253 10848 9259 10912
rect 9323 10848 9339 10912
rect 9403 10848 9419 10912
rect 9483 10848 9499 10912
rect 9563 10848 9569 10912
rect 9253 10847 9569 10848
rect 2038 10368 2354 10369
rect 2038 10304 2044 10368
rect 2108 10304 2124 10368
rect 2188 10304 2204 10368
rect 2268 10304 2284 10368
rect 2348 10304 2354 10368
rect 2038 10303 2354 10304
rect 4223 10368 4539 10369
rect 4223 10304 4229 10368
rect 4293 10304 4309 10368
rect 4373 10304 4389 10368
rect 4453 10304 4469 10368
rect 4533 10304 4539 10368
rect 4223 10303 4539 10304
rect 6408 10368 6724 10369
rect 6408 10304 6414 10368
rect 6478 10304 6494 10368
rect 6558 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6724 10368
rect 6408 10303 6724 10304
rect 8593 10368 8909 10369
rect 8593 10304 8599 10368
rect 8663 10304 8679 10368
rect 8743 10304 8759 10368
rect 8823 10304 8839 10368
rect 8903 10304 8909 10368
rect 8593 10303 8909 10304
rect 2698 9824 3014 9825
rect 2698 9760 2704 9824
rect 2768 9760 2784 9824
rect 2848 9760 2864 9824
rect 2928 9760 2944 9824
rect 3008 9760 3014 9824
rect 2698 9759 3014 9760
rect 4883 9824 5199 9825
rect 4883 9760 4889 9824
rect 4953 9760 4969 9824
rect 5033 9760 5049 9824
rect 5113 9760 5129 9824
rect 5193 9760 5199 9824
rect 4883 9759 5199 9760
rect 7068 9824 7384 9825
rect 7068 9760 7074 9824
rect 7138 9760 7154 9824
rect 7218 9760 7234 9824
rect 7298 9760 7314 9824
rect 7378 9760 7384 9824
rect 7068 9759 7384 9760
rect 9253 9824 9569 9825
rect 9253 9760 9259 9824
rect 9323 9760 9339 9824
rect 9403 9760 9419 9824
rect 9483 9760 9499 9824
rect 9563 9760 9569 9824
rect 9253 9759 9569 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 8017 9482 8083 9485
rect 8753 9482 8819 9485
rect 8017 9480 8819 9482
rect 8017 9424 8022 9480
rect 8078 9424 8758 9480
rect 8814 9424 8819 9480
rect 8017 9422 8819 9424
rect 8017 9419 8083 9422
rect 8753 9419 8819 9422
rect 2038 9280 2354 9281
rect 2038 9216 2044 9280
rect 2108 9216 2124 9280
rect 2188 9216 2204 9280
rect 2268 9216 2284 9280
rect 2348 9216 2354 9280
rect 2038 9215 2354 9216
rect 4223 9280 4539 9281
rect 4223 9216 4229 9280
rect 4293 9216 4309 9280
rect 4373 9216 4389 9280
rect 4453 9216 4469 9280
rect 4533 9216 4539 9280
rect 4223 9215 4539 9216
rect 6408 9280 6724 9281
rect 6408 9216 6414 9280
rect 6478 9216 6494 9280
rect 6558 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6724 9280
rect 6408 9215 6724 9216
rect 8593 9280 8909 9281
rect 8593 9216 8599 9280
rect 8663 9216 8679 9280
rect 8743 9216 8759 9280
rect 8823 9216 8839 9280
rect 8903 9216 8909 9280
rect 8593 9215 8909 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 0 8848 800 8878
rect 2698 8736 3014 8737
rect 2698 8672 2704 8736
rect 2768 8672 2784 8736
rect 2848 8672 2864 8736
rect 2928 8672 2944 8736
rect 3008 8672 3014 8736
rect 2698 8671 3014 8672
rect 4883 8736 5199 8737
rect 4883 8672 4889 8736
rect 4953 8672 4969 8736
rect 5033 8672 5049 8736
rect 5113 8672 5129 8736
rect 5193 8672 5199 8736
rect 4883 8671 5199 8672
rect 7068 8736 7384 8737
rect 7068 8672 7074 8736
rect 7138 8672 7154 8736
rect 7218 8672 7234 8736
rect 7298 8672 7314 8736
rect 7378 8672 7384 8736
rect 7068 8671 7384 8672
rect 9253 8736 9569 8737
rect 9253 8672 9259 8736
rect 9323 8672 9339 8736
rect 9403 8672 9419 8736
rect 9483 8672 9499 8736
rect 9563 8672 9569 8736
rect 9253 8671 9569 8672
rect 7097 8530 7163 8533
rect 8569 8530 8635 8533
rect 7097 8528 8635 8530
rect 7097 8472 7102 8528
rect 7158 8472 8574 8528
rect 8630 8472 8635 8528
rect 7097 8470 8635 8472
rect 7097 8467 7163 8470
rect 8569 8467 8635 8470
rect 9397 8258 9463 8261
rect 10164 8258 10964 8288
rect 9397 8256 10964 8258
rect 9397 8200 9402 8256
rect 9458 8200 10964 8256
rect 9397 8198 10964 8200
rect 9397 8195 9463 8198
rect 2038 8192 2354 8193
rect 2038 8128 2044 8192
rect 2108 8128 2124 8192
rect 2188 8128 2204 8192
rect 2268 8128 2284 8192
rect 2348 8128 2354 8192
rect 2038 8127 2354 8128
rect 4223 8192 4539 8193
rect 4223 8128 4229 8192
rect 4293 8128 4309 8192
rect 4373 8128 4389 8192
rect 4453 8128 4469 8192
rect 4533 8128 4539 8192
rect 4223 8127 4539 8128
rect 6408 8192 6724 8193
rect 6408 8128 6414 8192
rect 6478 8128 6494 8192
rect 6558 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6724 8192
rect 6408 8127 6724 8128
rect 8593 8192 8909 8193
rect 8593 8128 8599 8192
rect 8663 8128 8679 8192
rect 8743 8128 8759 8192
rect 8823 8128 8839 8192
rect 8903 8128 8909 8192
rect 10164 8168 10964 8198
rect 8593 8127 8909 8128
rect 7373 7986 7439 7989
rect 7649 7986 7715 7989
rect 9029 7986 9095 7989
rect 7373 7984 9095 7986
rect 7373 7928 7378 7984
rect 7434 7928 7654 7984
rect 7710 7928 9034 7984
rect 9090 7928 9095 7984
rect 7373 7926 9095 7928
rect 7373 7923 7439 7926
rect 7649 7923 7715 7926
rect 9029 7923 9095 7926
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 2698 7648 3014 7649
rect 2698 7584 2704 7648
rect 2768 7584 2784 7648
rect 2848 7584 2864 7648
rect 2928 7584 2944 7648
rect 3008 7584 3014 7648
rect 2698 7583 3014 7584
rect 4883 7648 5199 7649
rect 4883 7584 4889 7648
rect 4953 7584 4969 7648
rect 5033 7584 5049 7648
rect 5113 7584 5129 7648
rect 5193 7584 5199 7648
rect 4883 7583 5199 7584
rect 7068 7648 7384 7649
rect 7068 7584 7074 7648
rect 7138 7584 7154 7648
rect 7218 7584 7234 7648
rect 7298 7584 7314 7648
rect 7378 7584 7384 7648
rect 7068 7583 7384 7584
rect 9253 7648 9569 7649
rect 9253 7584 9259 7648
rect 9323 7584 9339 7648
rect 9403 7584 9419 7648
rect 9483 7584 9499 7648
rect 9563 7584 9569 7648
rect 9253 7583 9569 7584
rect 10164 7578 10964 7608
rect 9630 7518 10964 7578
rect 0 7488 800 7518
rect 7373 7442 7439 7445
rect 9630 7442 9690 7518
rect 10164 7488 10964 7518
rect 7373 7440 9690 7442
rect 7373 7384 7378 7440
rect 7434 7384 9690 7440
rect 7373 7382 9690 7384
rect 7373 7379 7439 7382
rect 2038 7104 2354 7105
rect 2038 7040 2044 7104
rect 2108 7040 2124 7104
rect 2188 7040 2204 7104
rect 2268 7040 2284 7104
rect 2348 7040 2354 7104
rect 2038 7039 2354 7040
rect 4223 7104 4539 7105
rect 4223 7040 4229 7104
rect 4293 7040 4309 7104
rect 4373 7040 4389 7104
rect 4453 7040 4469 7104
rect 4533 7040 4539 7104
rect 4223 7039 4539 7040
rect 6408 7104 6724 7105
rect 6408 7040 6414 7104
rect 6478 7040 6494 7104
rect 6558 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6724 7104
rect 6408 7039 6724 7040
rect 8593 7104 8909 7105
rect 8593 7040 8599 7104
rect 8663 7040 8679 7104
rect 8743 7040 8759 7104
rect 8823 7040 8839 7104
rect 8903 7040 8909 7104
rect 8593 7039 8909 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 9397 6898 9463 6901
rect 10164 6898 10964 6928
rect 9397 6896 10964 6898
rect 9397 6840 9402 6896
rect 9458 6840 10964 6896
rect 9397 6838 10964 6840
rect 9397 6835 9463 6838
rect 10164 6808 10964 6838
rect 2698 6560 3014 6561
rect 2698 6496 2704 6560
rect 2768 6496 2784 6560
rect 2848 6496 2864 6560
rect 2928 6496 2944 6560
rect 3008 6496 3014 6560
rect 2698 6495 3014 6496
rect 4883 6560 5199 6561
rect 4883 6496 4889 6560
rect 4953 6496 4969 6560
rect 5033 6496 5049 6560
rect 5113 6496 5129 6560
rect 5193 6496 5199 6560
rect 4883 6495 5199 6496
rect 7068 6560 7384 6561
rect 7068 6496 7074 6560
rect 7138 6496 7154 6560
rect 7218 6496 7234 6560
rect 7298 6496 7314 6560
rect 7378 6496 7384 6560
rect 7068 6495 7384 6496
rect 9253 6560 9569 6561
rect 9253 6496 9259 6560
rect 9323 6496 9339 6560
rect 9403 6496 9419 6560
rect 9483 6496 9499 6560
rect 9563 6496 9569 6560
rect 9253 6495 9569 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 7465 6218 7531 6221
rect 10164 6218 10964 6248
rect 7465 6216 10964 6218
rect 7465 6160 7470 6216
rect 7526 6160 10964 6216
rect 7465 6158 10964 6160
rect 0 6128 800 6158
rect 7465 6155 7531 6158
rect 10164 6128 10964 6158
rect 2038 6016 2354 6017
rect 2038 5952 2044 6016
rect 2108 5952 2124 6016
rect 2188 5952 2204 6016
rect 2268 5952 2284 6016
rect 2348 5952 2354 6016
rect 2038 5951 2354 5952
rect 4223 6016 4539 6017
rect 4223 5952 4229 6016
rect 4293 5952 4309 6016
rect 4373 5952 4389 6016
rect 4453 5952 4469 6016
rect 4533 5952 4539 6016
rect 4223 5951 4539 5952
rect 6408 6016 6724 6017
rect 6408 5952 6414 6016
rect 6478 5952 6494 6016
rect 6558 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6724 6016
rect 6408 5951 6724 5952
rect 8593 6016 8909 6017
rect 8593 5952 8599 6016
rect 8663 5952 8679 6016
rect 8743 5952 8759 6016
rect 8823 5952 8839 6016
rect 8903 5952 8909 6016
rect 8593 5951 8909 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 10164 5538 10964 5568
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 9630 5478 10964 5538
rect 2698 5472 3014 5473
rect 2698 5408 2704 5472
rect 2768 5408 2784 5472
rect 2848 5408 2864 5472
rect 2928 5408 2944 5472
rect 3008 5408 3014 5472
rect 2698 5407 3014 5408
rect 4883 5472 5199 5473
rect 4883 5408 4889 5472
rect 4953 5408 4969 5472
rect 5033 5408 5049 5472
rect 5113 5408 5129 5472
rect 5193 5408 5199 5472
rect 4883 5407 5199 5408
rect 7068 5472 7384 5473
rect 7068 5408 7074 5472
rect 7138 5408 7154 5472
rect 7218 5408 7234 5472
rect 7298 5408 7314 5472
rect 7378 5408 7384 5472
rect 7068 5407 7384 5408
rect 9253 5472 9569 5473
rect 9253 5408 9259 5472
rect 9323 5408 9339 5472
rect 9403 5408 9419 5472
rect 9483 5408 9499 5472
rect 9563 5408 9569 5472
rect 9253 5407 9569 5408
rect 2589 5266 2655 5269
rect 5257 5266 5323 5269
rect 2589 5264 5323 5266
rect 2589 5208 2594 5264
rect 2650 5208 5262 5264
rect 5318 5208 5323 5264
rect 2589 5206 5323 5208
rect 2589 5203 2655 5206
rect 5257 5203 5323 5206
rect 7189 5266 7255 5269
rect 9630 5266 9690 5478
rect 10164 5448 10964 5478
rect 7189 5264 9690 5266
rect 7189 5208 7194 5264
rect 7250 5208 9690 5264
rect 7189 5206 9690 5208
rect 7189 5203 7255 5206
rect 4521 5130 4587 5133
rect 4705 5130 4771 5133
rect 4521 5128 4771 5130
rect 4521 5072 4526 5128
rect 4582 5072 4710 5128
rect 4766 5072 4771 5128
rect 4521 5070 4771 5072
rect 4521 5067 4587 5070
rect 4705 5067 4771 5070
rect 2038 4928 2354 4929
rect 0 4858 800 4888
rect 2038 4864 2044 4928
rect 2108 4864 2124 4928
rect 2188 4864 2204 4928
rect 2268 4864 2284 4928
rect 2348 4864 2354 4928
rect 2038 4863 2354 4864
rect 4223 4928 4539 4929
rect 4223 4864 4229 4928
rect 4293 4864 4309 4928
rect 4373 4864 4389 4928
rect 4453 4864 4469 4928
rect 4533 4864 4539 4928
rect 4223 4863 4539 4864
rect 6408 4928 6724 4929
rect 6408 4864 6414 4928
rect 6478 4864 6494 4928
rect 6558 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6724 4928
rect 6408 4863 6724 4864
rect 8593 4928 8909 4929
rect 8593 4864 8599 4928
rect 8663 4864 8679 4928
rect 8743 4864 8759 4928
rect 8823 4864 8839 4928
rect 8903 4864 8909 4928
rect 8593 4863 8909 4864
rect 1209 4858 1275 4861
rect 0 4856 1275 4858
rect 0 4800 1214 4856
rect 1270 4800 1275 4856
rect 0 4798 1275 4800
rect 0 4768 800 4798
rect 1209 4795 1275 4798
rect 9581 4858 9647 4861
rect 10164 4858 10964 4888
rect 9581 4856 10964 4858
rect 9581 4800 9586 4856
rect 9642 4800 10964 4856
rect 9581 4798 10964 4800
rect 9581 4795 9647 4798
rect 10164 4768 10964 4798
rect 2698 4384 3014 4385
rect 2698 4320 2704 4384
rect 2768 4320 2784 4384
rect 2848 4320 2864 4384
rect 2928 4320 2944 4384
rect 3008 4320 3014 4384
rect 2698 4319 3014 4320
rect 4883 4384 5199 4385
rect 4883 4320 4889 4384
rect 4953 4320 4969 4384
rect 5033 4320 5049 4384
rect 5113 4320 5129 4384
rect 5193 4320 5199 4384
rect 4883 4319 5199 4320
rect 7068 4384 7384 4385
rect 7068 4320 7074 4384
rect 7138 4320 7154 4384
rect 7218 4320 7234 4384
rect 7298 4320 7314 4384
rect 7378 4320 7384 4384
rect 7068 4319 7384 4320
rect 9253 4384 9569 4385
rect 9253 4320 9259 4384
rect 9323 4320 9339 4384
rect 9403 4320 9419 4384
rect 9483 4320 9499 4384
rect 9563 4320 9569 4384
rect 9253 4319 9569 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 8293 4178 8359 4181
rect 10164 4178 10964 4208
rect 8293 4176 10964 4178
rect 8293 4120 8298 4176
rect 8354 4120 10964 4176
rect 8293 4118 10964 4120
rect 8293 4115 8359 4118
rect 10164 4088 10964 4118
rect 2038 3840 2354 3841
rect 2038 3776 2044 3840
rect 2108 3776 2124 3840
rect 2188 3776 2204 3840
rect 2268 3776 2284 3840
rect 2348 3776 2354 3840
rect 2038 3775 2354 3776
rect 4223 3840 4539 3841
rect 4223 3776 4229 3840
rect 4293 3776 4309 3840
rect 4373 3776 4389 3840
rect 4453 3776 4469 3840
rect 4533 3776 4539 3840
rect 4223 3775 4539 3776
rect 6408 3840 6724 3841
rect 6408 3776 6414 3840
rect 6478 3776 6494 3840
rect 6558 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6724 3840
rect 6408 3775 6724 3776
rect 8593 3840 8909 3841
rect 8593 3776 8599 3840
rect 8663 3776 8679 3840
rect 8743 3776 8759 3840
rect 8823 3776 8839 3840
rect 8903 3776 8909 3840
rect 8593 3775 8909 3776
rect 2698 3296 3014 3297
rect 2698 3232 2704 3296
rect 2768 3232 2784 3296
rect 2848 3232 2864 3296
rect 2928 3232 2944 3296
rect 3008 3232 3014 3296
rect 2698 3231 3014 3232
rect 4883 3296 5199 3297
rect 4883 3232 4889 3296
rect 4953 3232 4969 3296
rect 5033 3232 5049 3296
rect 5113 3232 5129 3296
rect 5193 3232 5199 3296
rect 4883 3231 5199 3232
rect 7068 3296 7384 3297
rect 7068 3232 7074 3296
rect 7138 3232 7154 3296
rect 7218 3232 7234 3296
rect 7298 3232 7314 3296
rect 7378 3232 7384 3296
rect 7068 3231 7384 3232
rect 9253 3296 9569 3297
rect 9253 3232 9259 3296
rect 9323 3232 9339 3296
rect 9403 3232 9419 3296
rect 9483 3232 9499 3296
rect 9563 3232 9569 3296
rect 9253 3231 9569 3232
rect 2038 2752 2354 2753
rect 2038 2688 2044 2752
rect 2108 2688 2124 2752
rect 2188 2688 2204 2752
rect 2268 2688 2284 2752
rect 2348 2688 2354 2752
rect 2038 2687 2354 2688
rect 4223 2752 4539 2753
rect 4223 2688 4229 2752
rect 4293 2688 4309 2752
rect 4373 2688 4389 2752
rect 4453 2688 4469 2752
rect 4533 2688 4539 2752
rect 4223 2687 4539 2688
rect 6408 2752 6724 2753
rect 6408 2688 6414 2752
rect 6478 2688 6494 2752
rect 6558 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6724 2752
rect 6408 2687 6724 2688
rect 8593 2752 8909 2753
rect 8593 2688 8599 2752
rect 8663 2688 8679 2752
rect 8743 2688 8759 2752
rect 8823 2688 8839 2752
rect 8903 2688 8909 2752
rect 8593 2687 8909 2688
rect 2698 2208 3014 2209
rect 2698 2144 2704 2208
rect 2768 2144 2784 2208
rect 2848 2144 2864 2208
rect 2928 2144 2944 2208
rect 3008 2144 3014 2208
rect 2698 2143 3014 2144
rect 4883 2208 5199 2209
rect 4883 2144 4889 2208
rect 4953 2144 4969 2208
rect 5033 2144 5049 2208
rect 5113 2144 5129 2208
rect 5193 2144 5199 2208
rect 4883 2143 5199 2144
rect 7068 2208 7384 2209
rect 7068 2144 7074 2208
rect 7138 2144 7154 2208
rect 7218 2144 7234 2208
rect 7298 2144 7314 2208
rect 7378 2144 7384 2208
rect 7068 2143 7384 2144
rect 9253 2208 9569 2209
rect 9253 2144 9259 2208
rect 9323 2144 9339 2208
rect 9403 2144 9419 2208
rect 9483 2144 9499 2208
rect 9563 2144 9569 2208
rect 9253 2143 9569 2144
<< via3 >>
rect 2704 10908 2768 10912
rect 2704 10852 2708 10908
rect 2708 10852 2764 10908
rect 2764 10852 2768 10908
rect 2704 10848 2768 10852
rect 2784 10908 2848 10912
rect 2784 10852 2788 10908
rect 2788 10852 2844 10908
rect 2844 10852 2848 10908
rect 2784 10848 2848 10852
rect 2864 10908 2928 10912
rect 2864 10852 2868 10908
rect 2868 10852 2924 10908
rect 2924 10852 2928 10908
rect 2864 10848 2928 10852
rect 2944 10908 3008 10912
rect 2944 10852 2948 10908
rect 2948 10852 3004 10908
rect 3004 10852 3008 10908
rect 2944 10848 3008 10852
rect 4889 10908 4953 10912
rect 4889 10852 4893 10908
rect 4893 10852 4949 10908
rect 4949 10852 4953 10908
rect 4889 10848 4953 10852
rect 4969 10908 5033 10912
rect 4969 10852 4973 10908
rect 4973 10852 5029 10908
rect 5029 10852 5033 10908
rect 4969 10848 5033 10852
rect 5049 10908 5113 10912
rect 5049 10852 5053 10908
rect 5053 10852 5109 10908
rect 5109 10852 5113 10908
rect 5049 10848 5113 10852
rect 5129 10908 5193 10912
rect 5129 10852 5133 10908
rect 5133 10852 5189 10908
rect 5189 10852 5193 10908
rect 5129 10848 5193 10852
rect 7074 10908 7138 10912
rect 7074 10852 7078 10908
rect 7078 10852 7134 10908
rect 7134 10852 7138 10908
rect 7074 10848 7138 10852
rect 7154 10908 7218 10912
rect 7154 10852 7158 10908
rect 7158 10852 7214 10908
rect 7214 10852 7218 10908
rect 7154 10848 7218 10852
rect 7234 10908 7298 10912
rect 7234 10852 7238 10908
rect 7238 10852 7294 10908
rect 7294 10852 7298 10908
rect 7234 10848 7298 10852
rect 7314 10908 7378 10912
rect 7314 10852 7318 10908
rect 7318 10852 7374 10908
rect 7374 10852 7378 10908
rect 7314 10848 7378 10852
rect 9259 10908 9323 10912
rect 9259 10852 9263 10908
rect 9263 10852 9319 10908
rect 9319 10852 9323 10908
rect 9259 10848 9323 10852
rect 9339 10908 9403 10912
rect 9339 10852 9343 10908
rect 9343 10852 9399 10908
rect 9399 10852 9403 10908
rect 9339 10848 9403 10852
rect 9419 10908 9483 10912
rect 9419 10852 9423 10908
rect 9423 10852 9479 10908
rect 9479 10852 9483 10908
rect 9419 10848 9483 10852
rect 9499 10908 9563 10912
rect 9499 10852 9503 10908
rect 9503 10852 9559 10908
rect 9559 10852 9563 10908
rect 9499 10848 9563 10852
rect 2044 10364 2108 10368
rect 2044 10308 2048 10364
rect 2048 10308 2104 10364
rect 2104 10308 2108 10364
rect 2044 10304 2108 10308
rect 2124 10364 2188 10368
rect 2124 10308 2128 10364
rect 2128 10308 2184 10364
rect 2184 10308 2188 10364
rect 2124 10304 2188 10308
rect 2204 10364 2268 10368
rect 2204 10308 2208 10364
rect 2208 10308 2264 10364
rect 2264 10308 2268 10364
rect 2204 10304 2268 10308
rect 2284 10364 2348 10368
rect 2284 10308 2288 10364
rect 2288 10308 2344 10364
rect 2344 10308 2348 10364
rect 2284 10304 2348 10308
rect 4229 10364 4293 10368
rect 4229 10308 4233 10364
rect 4233 10308 4289 10364
rect 4289 10308 4293 10364
rect 4229 10304 4293 10308
rect 4309 10364 4373 10368
rect 4309 10308 4313 10364
rect 4313 10308 4369 10364
rect 4369 10308 4373 10364
rect 4309 10304 4373 10308
rect 4389 10364 4453 10368
rect 4389 10308 4393 10364
rect 4393 10308 4449 10364
rect 4449 10308 4453 10364
rect 4389 10304 4453 10308
rect 4469 10364 4533 10368
rect 4469 10308 4473 10364
rect 4473 10308 4529 10364
rect 4529 10308 4533 10364
rect 4469 10304 4533 10308
rect 6414 10364 6478 10368
rect 6414 10308 6418 10364
rect 6418 10308 6474 10364
rect 6474 10308 6478 10364
rect 6414 10304 6478 10308
rect 6494 10364 6558 10368
rect 6494 10308 6498 10364
rect 6498 10308 6554 10364
rect 6554 10308 6558 10364
rect 6494 10304 6558 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 8599 10364 8663 10368
rect 8599 10308 8603 10364
rect 8603 10308 8659 10364
rect 8659 10308 8663 10364
rect 8599 10304 8663 10308
rect 8679 10364 8743 10368
rect 8679 10308 8683 10364
rect 8683 10308 8739 10364
rect 8739 10308 8743 10364
rect 8679 10304 8743 10308
rect 8759 10364 8823 10368
rect 8759 10308 8763 10364
rect 8763 10308 8819 10364
rect 8819 10308 8823 10364
rect 8759 10304 8823 10308
rect 8839 10364 8903 10368
rect 8839 10308 8843 10364
rect 8843 10308 8899 10364
rect 8899 10308 8903 10364
rect 8839 10304 8903 10308
rect 2704 9820 2768 9824
rect 2704 9764 2708 9820
rect 2708 9764 2764 9820
rect 2764 9764 2768 9820
rect 2704 9760 2768 9764
rect 2784 9820 2848 9824
rect 2784 9764 2788 9820
rect 2788 9764 2844 9820
rect 2844 9764 2848 9820
rect 2784 9760 2848 9764
rect 2864 9820 2928 9824
rect 2864 9764 2868 9820
rect 2868 9764 2924 9820
rect 2924 9764 2928 9820
rect 2864 9760 2928 9764
rect 2944 9820 3008 9824
rect 2944 9764 2948 9820
rect 2948 9764 3004 9820
rect 3004 9764 3008 9820
rect 2944 9760 3008 9764
rect 4889 9820 4953 9824
rect 4889 9764 4893 9820
rect 4893 9764 4949 9820
rect 4949 9764 4953 9820
rect 4889 9760 4953 9764
rect 4969 9820 5033 9824
rect 4969 9764 4973 9820
rect 4973 9764 5029 9820
rect 5029 9764 5033 9820
rect 4969 9760 5033 9764
rect 5049 9820 5113 9824
rect 5049 9764 5053 9820
rect 5053 9764 5109 9820
rect 5109 9764 5113 9820
rect 5049 9760 5113 9764
rect 5129 9820 5193 9824
rect 5129 9764 5133 9820
rect 5133 9764 5189 9820
rect 5189 9764 5193 9820
rect 5129 9760 5193 9764
rect 7074 9820 7138 9824
rect 7074 9764 7078 9820
rect 7078 9764 7134 9820
rect 7134 9764 7138 9820
rect 7074 9760 7138 9764
rect 7154 9820 7218 9824
rect 7154 9764 7158 9820
rect 7158 9764 7214 9820
rect 7214 9764 7218 9820
rect 7154 9760 7218 9764
rect 7234 9820 7298 9824
rect 7234 9764 7238 9820
rect 7238 9764 7294 9820
rect 7294 9764 7298 9820
rect 7234 9760 7298 9764
rect 7314 9820 7378 9824
rect 7314 9764 7318 9820
rect 7318 9764 7374 9820
rect 7374 9764 7378 9820
rect 7314 9760 7378 9764
rect 9259 9820 9323 9824
rect 9259 9764 9263 9820
rect 9263 9764 9319 9820
rect 9319 9764 9323 9820
rect 9259 9760 9323 9764
rect 9339 9820 9403 9824
rect 9339 9764 9343 9820
rect 9343 9764 9399 9820
rect 9399 9764 9403 9820
rect 9339 9760 9403 9764
rect 9419 9820 9483 9824
rect 9419 9764 9423 9820
rect 9423 9764 9479 9820
rect 9479 9764 9483 9820
rect 9419 9760 9483 9764
rect 9499 9820 9563 9824
rect 9499 9764 9503 9820
rect 9503 9764 9559 9820
rect 9559 9764 9563 9820
rect 9499 9760 9563 9764
rect 2044 9276 2108 9280
rect 2044 9220 2048 9276
rect 2048 9220 2104 9276
rect 2104 9220 2108 9276
rect 2044 9216 2108 9220
rect 2124 9276 2188 9280
rect 2124 9220 2128 9276
rect 2128 9220 2184 9276
rect 2184 9220 2188 9276
rect 2124 9216 2188 9220
rect 2204 9276 2268 9280
rect 2204 9220 2208 9276
rect 2208 9220 2264 9276
rect 2264 9220 2268 9276
rect 2204 9216 2268 9220
rect 2284 9276 2348 9280
rect 2284 9220 2288 9276
rect 2288 9220 2344 9276
rect 2344 9220 2348 9276
rect 2284 9216 2348 9220
rect 4229 9276 4293 9280
rect 4229 9220 4233 9276
rect 4233 9220 4289 9276
rect 4289 9220 4293 9276
rect 4229 9216 4293 9220
rect 4309 9276 4373 9280
rect 4309 9220 4313 9276
rect 4313 9220 4369 9276
rect 4369 9220 4373 9276
rect 4309 9216 4373 9220
rect 4389 9276 4453 9280
rect 4389 9220 4393 9276
rect 4393 9220 4449 9276
rect 4449 9220 4453 9276
rect 4389 9216 4453 9220
rect 4469 9276 4533 9280
rect 4469 9220 4473 9276
rect 4473 9220 4529 9276
rect 4529 9220 4533 9276
rect 4469 9216 4533 9220
rect 6414 9276 6478 9280
rect 6414 9220 6418 9276
rect 6418 9220 6474 9276
rect 6474 9220 6478 9276
rect 6414 9216 6478 9220
rect 6494 9276 6558 9280
rect 6494 9220 6498 9276
rect 6498 9220 6554 9276
rect 6554 9220 6558 9276
rect 6494 9216 6558 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 8599 9276 8663 9280
rect 8599 9220 8603 9276
rect 8603 9220 8659 9276
rect 8659 9220 8663 9276
rect 8599 9216 8663 9220
rect 8679 9276 8743 9280
rect 8679 9220 8683 9276
rect 8683 9220 8739 9276
rect 8739 9220 8743 9276
rect 8679 9216 8743 9220
rect 8759 9276 8823 9280
rect 8759 9220 8763 9276
rect 8763 9220 8819 9276
rect 8819 9220 8823 9276
rect 8759 9216 8823 9220
rect 8839 9276 8903 9280
rect 8839 9220 8843 9276
rect 8843 9220 8899 9276
rect 8899 9220 8903 9276
rect 8839 9216 8903 9220
rect 2704 8732 2768 8736
rect 2704 8676 2708 8732
rect 2708 8676 2764 8732
rect 2764 8676 2768 8732
rect 2704 8672 2768 8676
rect 2784 8732 2848 8736
rect 2784 8676 2788 8732
rect 2788 8676 2844 8732
rect 2844 8676 2848 8732
rect 2784 8672 2848 8676
rect 2864 8732 2928 8736
rect 2864 8676 2868 8732
rect 2868 8676 2924 8732
rect 2924 8676 2928 8732
rect 2864 8672 2928 8676
rect 2944 8732 3008 8736
rect 2944 8676 2948 8732
rect 2948 8676 3004 8732
rect 3004 8676 3008 8732
rect 2944 8672 3008 8676
rect 4889 8732 4953 8736
rect 4889 8676 4893 8732
rect 4893 8676 4949 8732
rect 4949 8676 4953 8732
rect 4889 8672 4953 8676
rect 4969 8732 5033 8736
rect 4969 8676 4973 8732
rect 4973 8676 5029 8732
rect 5029 8676 5033 8732
rect 4969 8672 5033 8676
rect 5049 8732 5113 8736
rect 5049 8676 5053 8732
rect 5053 8676 5109 8732
rect 5109 8676 5113 8732
rect 5049 8672 5113 8676
rect 5129 8732 5193 8736
rect 5129 8676 5133 8732
rect 5133 8676 5189 8732
rect 5189 8676 5193 8732
rect 5129 8672 5193 8676
rect 7074 8732 7138 8736
rect 7074 8676 7078 8732
rect 7078 8676 7134 8732
rect 7134 8676 7138 8732
rect 7074 8672 7138 8676
rect 7154 8732 7218 8736
rect 7154 8676 7158 8732
rect 7158 8676 7214 8732
rect 7214 8676 7218 8732
rect 7154 8672 7218 8676
rect 7234 8732 7298 8736
rect 7234 8676 7238 8732
rect 7238 8676 7294 8732
rect 7294 8676 7298 8732
rect 7234 8672 7298 8676
rect 7314 8732 7378 8736
rect 7314 8676 7318 8732
rect 7318 8676 7374 8732
rect 7374 8676 7378 8732
rect 7314 8672 7378 8676
rect 9259 8732 9323 8736
rect 9259 8676 9263 8732
rect 9263 8676 9319 8732
rect 9319 8676 9323 8732
rect 9259 8672 9323 8676
rect 9339 8732 9403 8736
rect 9339 8676 9343 8732
rect 9343 8676 9399 8732
rect 9399 8676 9403 8732
rect 9339 8672 9403 8676
rect 9419 8732 9483 8736
rect 9419 8676 9423 8732
rect 9423 8676 9479 8732
rect 9479 8676 9483 8732
rect 9419 8672 9483 8676
rect 9499 8732 9563 8736
rect 9499 8676 9503 8732
rect 9503 8676 9559 8732
rect 9559 8676 9563 8732
rect 9499 8672 9563 8676
rect 2044 8188 2108 8192
rect 2044 8132 2048 8188
rect 2048 8132 2104 8188
rect 2104 8132 2108 8188
rect 2044 8128 2108 8132
rect 2124 8188 2188 8192
rect 2124 8132 2128 8188
rect 2128 8132 2184 8188
rect 2184 8132 2188 8188
rect 2124 8128 2188 8132
rect 2204 8188 2268 8192
rect 2204 8132 2208 8188
rect 2208 8132 2264 8188
rect 2264 8132 2268 8188
rect 2204 8128 2268 8132
rect 2284 8188 2348 8192
rect 2284 8132 2288 8188
rect 2288 8132 2344 8188
rect 2344 8132 2348 8188
rect 2284 8128 2348 8132
rect 4229 8188 4293 8192
rect 4229 8132 4233 8188
rect 4233 8132 4289 8188
rect 4289 8132 4293 8188
rect 4229 8128 4293 8132
rect 4309 8188 4373 8192
rect 4309 8132 4313 8188
rect 4313 8132 4369 8188
rect 4369 8132 4373 8188
rect 4309 8128 4373 8132
rect 4389 8188 4453 8192
rect 4389 8132 4393 8188
rect 4393 8132 4449 8188
rect 4449 8132 4453 8188
rect 4389 8128 4453 8132
rect 4469 8188 4533 8192
rect 4469 8132 4473 8188
rect 4473 8132 4529 8188
rect 4529 8132 4533 8188
rect 4469 8128 4533 8132
rect 6414 8188 6478 8192
rect 6414 8132 6418 8188
rect 6418 8132 6474 8188
rect 6474 8132 6478 8188
rect 6414 8128 6478 8132
rect 6494 8188 6558 8192
rect 6494 8132 6498 8188
rect 6498 8132 6554 8188
rect 6554 8132 6558 8188
rect 6494 8128 6558 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 8599 8188 8663 8192
rect 8599 8132 8603 8188
rect 8603 8132 8659 8188
rect 8659 8132 8663 8188
rect 8599 8128 8663 8132
rect 8679 8188 8743 8192
rect 8679 8132 8683 8188
rect 8683 8132 8739 8188
rect 8739 8132 8743 8188
rect 8679 8128 8743 8132
rect 8759 8188 8823 8192
rect 8759 8132 8763 8188
rect 8763 8132 8819 8188
rect 8819 8132 8823 8188
rect 8759 8128 8823 8132
rect 8839 8188 8903 8192
rect 8839 8132 8843 8188
rect 8843 8132 8899 8188
rect 8899 8132 8903 8188
rect 8839 8128 8903 8132
rect 2704 7644 2768 7648
rect 2704 7588 2708 7644
rect 2708 7588 2764 7644
rect 2764 7588 2768 7644
rect 2704 7584 2768 7588
rect 2784 7644 2848 7648
rect 2784 7588 2788 7644
rect 2788 7588 2844 7644
rect 2844 7588 2848 7644
rect 2784 7584 2848 7588
rect 2864 7644 2928 7648
rect 2864 7588 2868 7644
rect 2868 7588 2924 7644
rect 2924 7588 2928 7644
rect 2864 7584 2928 7588
rect 2944 7644 3008 7648
rect 2944 7588 2948 7644
rect 2948 7588 3004 7644
rect 3004 7588 3008 7644
rect 2944 7584 3008 7588
rect 4889 7644 4953 7648
rect 4889 7588 4893 7644
rect 4893 7588 4949 7644
rect 4949 7588 4953 7644
rect 4889 7584 4953 7588
rect 4969 7644 5033 7648
rect 4969 7588 4973 7644
rect 4973 7588 5029 7644
rect 5029 7588 5033 7644
rect 4969 7584 5033 7588
rect 5049 7644 5113 7648
rect 5049 7588 5053 7644
rect 5053 7588 5109 7644
rect 5109 7588 5113 7644
rect 5049 7584 5113 7588
rect 5129 7644 5193 7648
rect 5129 7588 5133 7644
rect 5133 7588 5189 7644
rect 5189 7588 5193 7644
rect 5129 7584 5193 7588
rect 7074 7644 7138 7648
rect 7074 7588 7078 7644
rect 7078 7588 7134 7644
rect 7134 7588 7138 7644
rect 7074 7584 7138 7588
rect 7154 7644 7218 7648
rect 7154 7588 7158 7644
rect 7158 7588 7214 7644
rect 7214 7588 7218 7644
rect 7154 7584 7218 7588
rect 7234 7644 7298 7648
rect 7234 7588 7238 7644
rect 7238 7588 7294 7644
rect 7294 7588 7298 7644
rect 7234 7584 7298 7588
rect 7314 7644 7378 7648
rect 7314 7588 7318 7644
rect 7318 7588 7374 7644
rect 7374 7588 7378 7644
rect 7314 7584 7378 7588
rect 9259 7644 9323 7648
rect 9259 7588 9263 7644
rect 9263 7588 9319 7644
rect 9319 7588 9323 7644
rect 9259 7584 9323 7588
rect 9339 7644 9403 7648
rect 9339 7588 9343 7644
rect 9343 7588 9399 7644
rect 9399 7588 9403 7644
rect 9339 7584 9403 7588
rect 9419 7644 9483 7648
rect 9419 7588 9423 7644
rect 9423 7588 9479 7644
rect 9479 7588 9483 7644
rect 9419 7584 9483 7588
rect 9499 7644 9563 7648
rect 9499 7588 9503 7644
rect 9503 7588 9559 7644
rect 9559 7588 9563 7644
rect 9499 7584 9563 7588
rect 2044 7100 2108 7104
rect 2044 7044 2048 7100
rect 2048 7044 2104 7100
rect 2104 7044 2108 7100
rect 2044 7040 2108 7044
rect 2124 7100 2188 7104
rect 2124 7044 2128 7100
rect 2128 7044 2184 7100
rect 2184 7044 2188 7100
rect 2124 7040 2188 7044
rect 2204 7100 2268 7104
rect 2204 7044 2208 7100
rect 2208 7044 2264 7100
rect 2264 7044 2268 7100
rect 2204 7040 2268 7044
rect 2284 7100 2348 7104
rect 2284 7044 2288 7100
rect 2288 7044 2344 7100
rect 2344 7044 2348 7100
rect 2284 7040 2348 7044
rect 4229 7100 4293 7104
rect 4229 7044 4233 7100
rect 4233 7044 4289 7100
rect 4289 7044 4293 7100
rect 4229 7040 4293 7044
rect 4309 7100 4373 7104
rect 4309 7044 4313 7100
rect 4313 7044 4369 7100
rect 4369 7044 4373 7100
rect 4309 7040 4373 7044
rect 4389 7100 4453 7104
rect 4389 7044 4393 7100
rect 4393 7044 4449 7100
rect 4449 7044 4453 7100
rect 4389 7040 4453 7044
rect 4469 7100 4533 7104
rect 4469 7044 4473 7100
rect 4473 7044 4529 7100
rect 4529 7044 4533 7100
rect 4469 7040 4533 7044
rect 6414 7100 6478 7104
rect 6414 7044 6418 7100
rect 6418 7044 6474 7100
rect 6474 7044 6478 7100
rect 6414 7040 6478 7044
rect 6494 7100 6558 7104
rect 6494 7044 6498 7100
rect 6498 7044 6554 7100
rect 6554 7044 6558 7100
rect 6494 7040 6558 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 8599 7100 8663 7104
rect 8599 7044 8603 7100
rect 8603 7044 8659 7100
rect 8659 7044 8663 7100
rect 8599 7040 8663 7044
rect 8679 7100 8743 7104
rect 8679 7044 8683 7100
rect 8683 7044 8739 7100
rect 8739 7044 8743 7100
rect 8679 7040 8743 7044
rect 8759 7100 8823 7104
rect 8759 7044 8763 7100
rect 8763 7044 8819 7100
rect 8819 7044 8823 7100
rect 8759 7040 8823 7044
rect 8839 7100 8903 7104
rect 8839 7044 8843 7100
rect 8843 7044 8899 7100
rect 8899 7044 8903 7100
rect 8839 7040 8903 7044
rect 2704 6556 2768 6560
rect 2704 6500 2708 6556
rect 2708 6500 2764 6556
rect 2764 6500 2768 6556
rect 2704 6496 2768 6500
rect 2784 6556 2848 6560
rect 2784 6500 2788 6556
rect 2788 6500 2844 6556
rect 2844 6500 2848 6556
rect 2784 6496 2848 6500
rect 2864 6556 2928 6560
rect 2864 6500 2868 6556
rect 2868 6500 2924 6556
rect 2924 6500 2928 6556
rect 2864 6496 2928 6500
rect 2944 6556 3008 6560
rect 2944 6500 2948 6556
rect 2948 6500 3004 6556
rect 3004 6500 3008 6556
rect 2944 6496 3008 6500
rect 4889 6556 4953 6560
rect 4889 6500 4893 6556
rect 4893 6500 4949 6556
rect 4949 6500 4953 6556
rect 4889 6496 4953 6500
rect 4969 6556 5033 6560
rect 4969 6500 4973 6556
rect 4973 6500 5029 6556
rect 5029 6500 5033 6556
rect 4969 6496 5033 6500
rect 5049 6556 5113 6560
rect 5049 6500 5053 6556
rect 5053 6500 5109 6556
rect 5109 6500 5113 6556
rect 5049 6496 5113 6500
rect 5129 6556 5193 6560
rect 5129 6500 5133 6556
rect 5133 6500 5189 6556
rect 5189 6500 5193 6556
rect 5129 6496 5193 6500
rect 7074 6556 7138 6560
rect 7074 6500 7078 6556
rect 7078 6500 7134 6556
rect 7134 6500 7138 6556
rect 7074 6496 7138 6500
rect 7154 6556 7218 6560
rect 7154 6500 7158 6556
rect 7158 6500 7214 6556
rect 7214 6500 7218 6556
rect 7154 6496 7218 6500
rect 7234 6556 7298 6560
rect 7234 6500 7238 6556
rect 7238 6500 7294 6556
rect 7294 6500 7298 6556
rect 7234 6496 7298 6500
rect 7314 6556 7378 6560
rect 7314 6500 7318 6556
rect 7318 6500 7374 6556
rect 7374 6500 7378 6556
rect 7314 6496 7378 6500
rect 9259 6556 9323 6560
rect 9259 6500 9263 6556
rect 9263 6500 9319 6556
rect 9319 6500 9323 6556
rect 9259 6496 9323 6500
rect 9339 6556 9403 6560
rect 9339 6500 9343 6556
rect 9343 6500 9399 6556
rect 9399 6500 9403 6556
rect 9339 6496 9403 6500
rect 9419 6556 9483 6560
rect 9419 6500 9423 6556
rect 9423 6500 9479 6556
rect 9479 6500 9483 6556
rect 9419 6496 9483 6500
rect 9499 6556 9563 6560
rect 9499 6500 9503 6556
rect 9503 6500 9559 6556
rect 9559 6500 9563 6556
rect 9499 6496 9563 6500
rect 2044 6012 2108 6016
rect 2044 5956 2048 6012
rect 2048 5956 2104 6012
rect 2104 5956 2108 6012
rect 2044 5952 2108 5956
rect 2124 6012 2188 6016
rect 2124 5956 2128 6012
rect 2128 5956 2184 6012
rect 2184 5956 2188 6012
rect 2124 5952 2188 5956
rect 2204 6012 2268 6016
rect 2204 5956 2208 6012
rect 2208 5956 2264 6012
rect 2264 5956 2268 6012
rect 2204 5952 2268 5956
rect 2284 6012 2348 6016
rect 2284 5956 2288 6012
rect 2288 5956 2344 6012
rect 2344 5956 2348 6012
rect 2284 5952 2348 5956
rect 4229 6012 4293 6016
rect 4229 5956 4233 6012
rect 4233 5956 4289 6012
rect 4289 5956 4293 6012
rect 4229 5952 4293 5956
rect 4309 6012 4373 6016
rect 4309 5956 4313 6012
rect 4313 5956 4369 6012
rect 4369 5956 4373 6012
rect 4309 5952 4373 5956
rect 4389 6012 4453 6016
rect 4389 5956 4393 6012
rect 4393 5956 4449 6012
rect 4449 5956 4453 6012
rect 4389 5952 4453 5956
rect 4469 6012 4533 6016
rect 4469 5956 4473 6012
rect 4473 5956 4529 6012
rect 4529 5956 4533 6012
rect 4469 5952 4533 5956
rect 6414 6012 6478 6016
rect 6414 5956 6418 6012
rect 6418 5956 6474 6012
rect 6474 5956 6478 6012
rect 6414 5952 6478 5956
rect 6494 6012 6558 6016
rect 6494 5956 6498 6012
rect 6498 5956 6554 6012
rect 6554 5956 6558 6012
rect 6494 5952 6558 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 8599 6012 8663 6016
rect 8599 5956 8603 6012
rect 8603 5956 8659 6012
rect 8659 5956 8663 6012
rect 8599 5952 8663 5956
rect 8679 6012 8743 6016
rect 8679 5956 8683 6012
rect 8683 5956 8739 6012
rect 8739 5956 8743 6012
rect 8679 5952 8743 5956
rect 8759 6012 8823 6016
rect 8759 5956 8763 6012
rect 8763 5956 8819 6012
rect 8819 5956 8823 6012
rect 8759 5952 8823 5956
rect 8839 6012 8903 6016
rect 8839 5956 8843 6012
rect 8843 5956 8899 6012
rect 8899 5956 8903 6012
rect 8839 5952 8903 5956
rect 2704 5468 2768 5472
rect 2704 5412 2708 5468
rect 2708 5412 2764 5468
rect 2764 5412 2768 5468
rect 2704 5408 2768 5412
rect 2784 5468 2848 5472
rect 2784 5412 2788 5468
rect 2788 5412 2844 5468
rect 2844 5412 2848 5468
rect 2784 5408 2848 5412
rect 2864 5468 2928 5472
rect 2864 5412 2868 5468
rect 2868 5412 2924 5468
rect 2924 5412 2928 5468
rect 2864 5408 2928 5412
rect 2944 5468 3008 5472
rect 2944 5412 2948 5468
rect 2948 5412 3004 5468
rect 3004 5412 3008 5468
rect 2944 5408 3008 5412
rect 4889 5468 4953 5472
rect 4889 5412 4893 5468
rect 4893 5412 4949 5468
rect 4949 5412 4953 5468
rect 4889 5408 4953 5412
rect 4969 5468 5033 5472
rect 4969 5412 4973 5468
rect 4973 5412 5029 5468
rect 5029 5412 5033 5468
rect 4969 5408 5033 5412
rect 5049 5468 5113 5472
rect 5049 5412 5053 5468
rect 5053 5412 5109 5468
rect 5109 5412 5113 5468
rect 5049 5408 5113 5412
rect 5129 5468 5193 5472
rect 5129 5412 5133 5468
rect 5133 5412 5189 5468
rect 5189 5412 5193 5468
rect 5129 5408 5193 5412
rect 7074 5468 7138 5472
rect 7074 5412 7078 5468
rect 7078 5412 7134 5468
rect 7134 5412 7138 5468
rect 7074 5408 7138 5412
rect 7154 5468 7218 5472
rect 7154 5412 7158 5468
rect 7158 5412 7214 5468
rect 7214 5412 7218 5468
rect 7154 5408 7218 5412
rect 7234 5468 7298 5472
rect 7234 5412 7238 5468
rect 7238 5412 7294 5468
rect 7294 5412 7298 5468
rect 7234 5408 7298 5412
rect 7314 5468 7378 5472
rect 7314 5412 7318 5468
rect 7318 5412 7374 5468
rect 7374 5412 7378 5468
rect 7314 5408 7378 5412
rect 9259 5468 9323 5472
rect 9259 5412 9263 5468
rect 9263 5412 9319 5468
rect 9319 5412 9323 5468
rect 9259 5408 9323 5412
rect 9339 5468 9403 5472
rect 9339 5412 9343 5468
rect 9343 5412 9399 5468
rect 9399 5412 9403 5468
rect 9339 5408 9403 5412
rect 9419 5468 9483 5472
rect 9419 5412 9423 5468
rect 9423 5412 9479 5468
rect 9479 5412 9483 5468
rect 9419 5408 9483 5412
rect 9499 5468 9563 5472
rect 9499 5412 9503 5468
rect 9503 5412 9559 5468
rect 9559 5412 9563 5468
rect 9499 5408 9563 5412
rect 2044 4924 2108 4928
rect 2044 4868 2048 4924
rect 2048 4868 2104 4924
rect 2104 4868 2108 4924
rect 2044 4864 2108 4868
rect 2124 4924 2188 4928
rect 2124 4868 2128 4924
rect 2128 4868 2184 4924
rect 2184 4868 2188 4924
rect 2124 4864 2188 4868
rect 2204 4924 2268 4928
rect 2204 4868 2208 4924
rect 2208 4868 2264 4924
rect 2264 4868 2268 4924
rect 2204 4864 2268 4868
rect 2284 4924 2348 4928
rect 2284 4868 2288 4924
rect 2288 4868 2344 4924
rect 2344 4868 2348 4924
rect 2284 4864 2348 4868
rect 4229 4924 4293 4928
rect 4229 4868 4233 4924
rect 4233 4868 4289 4924
rect 4289 4868 4293 4924
rect 4229 4864 4293 4868
rect 4309 4924 4373 4928
rect 4309 4868 4313 4924
rect 4313 4868 4369 4924
rect 4369 4868 4373 4924
rect 4309 4864 4373 4868
rect 4389 4924 4453 4928
rect 4389 4868 4393 4924
rect 4393 4868 4449 4924
rect 4449 4868 4453 4924
rect 4389 4864 4453 4868
rect 4469 4924 4533 4928
rect 4469 4868 4473 4924
rect 4473 4868 4529 4924
rect 4529 4868 4533 4924
rect 4469 4864 4533 4868
rect 6414 4924 6478 4928
rect 6414 4868 6418 4924
rect 6418 4868 6474 4924
rect 6474 4868 6478 4924
rect 6414 4864 6478 4868
rect 6494 4924 6558 4928
rect 6494 4868 6498 4924
rect 6498 4868 6554 4924
rect 6554 4868 6558 4924
rect 6494 4864 6558 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 8599 4924 8663 4928
rect 8599 4868 8603 4924
rect 8603 4868 8659 4924
rect 8659 4868 8663 4924
rect 8599 4864 8663 4868
rect 8679 4924 8743 4928
rect 8679 4868 8683 4924
rect 8683 4868 8739 4924
rect 8739 4868 8743 4924
rect 8679 4864 8743 4868
rect 8759 4924 8823 4928
rect 8759 4868 8763 4924
rect 8763 4868 8819 4924
rect 8819 4868 8823 4924
rect 8759 4864 8823 4868
rect 8839 4924 8903 4928
rect 8839 4868 8843 4924
rect 8843 4868 8899 4924
rect 8899 4868 8903 4924
rect 8839 4864 8903 4868
rect 2704 4380 2768 4384
rect 2704 4324 2708 4380
rect 2708 4324 2764 4380
rect 2764 4324 2768 4380
rect 2704 4320 2768 4324
rect 2784 4380 2848 4384
rect 2784 4324 2788 4380
rect 2788 4324 2844 4380
rect 2844 4324 2848 4380
rect 2784 4320 2848 4324
rect 2864 4380 2928 4384
rect 2864 4324 2868 4380
rect 2868 4324 2924 4380
rect 2924 4324 2928 4380
rect 2864 4320 2928 4324
rect 2944 4380 3008 4384
rect 2944 4324 2948 4380
rect 2948 4324 3004 4380
rect 3004 4324 3008 4380
rect 2944 4320 3008 4324
rect 4889 4380 4953 4384
rect 4889 4324 4893 4380
rect 4893 4324 4949 4380
rect 4949 4324 4953 4380
rect 4889 4320 4953 4324
rect 4969 4380 5033 4384
rect 4969 4324 4973 4380
rect 4973 4324 5029 4380
rect 5029 4324 5033 4380
rect 4969 4320 5033 4324
rect 5049 4380 5113 4384
rect 5049 4324 5053 4380
rect 5053 4324 5109 4380
rect 5109 4324 5113 4380
rect 5049 4320 5113 4324
rect 5129 4380 5193 4384
rect 5129 4324 5133 4380
rect 5133 4324 5189 4380
rect 5189 4324 5193 4380
rect 5129 4320 5193 4324
rect 7074 4380 7138 4384
rect 7074 4324 7078 4380
rect 7078 4324 7134 4380
rect 7134 4324 7138 4380
rect 7074 4320 7138 4324
rect 7154 4380 7218 4384
rect 7154 4324 7158 4380
rect 7158 4324 7214 4380
rect 7214 4324 7218 4380
rect 7154 4320 7218 4324
rect 7234 4380 7298 4384
rect 7234 4324 7238 4380
rect 7238 4324 7294 4380
rect 7294 4324 7298 4380
rect 7234 4320 7298 4324
rect 7314 4380 7378 4384
rect 7314 4324 7318 4380
rect 7318 4324 7374 4380
rect 7374 4324 7378 4380
rect 7314 4320 7378 4324
rect 9259 4380 9323 4384
rect 9259 4324 9263 4380
rect 9263 4324 9319 4380
rect 9319 4324 9323 4380
rect 9259 4320 9323 4324
rect 9339 4380 9403 4384
rect 9339 4324 9343 4380
rect 9343 4324 9399 4380
rect 9399 4324 9403 4380
rect 9339 4320 9403 4324
rect 9419 4380 9483 4384
rect 9419 4324 9423 4380
rect 9423 4324 9479 4380
rect 9479 4324 9483 4380
rect 9419 4320 9483 4324
rect 9499 4380 9563 4384
rect 9499 4324 9503 4380
rect 9503 4324 9559 4380
rect 9559 4324 9563 4380
rect 9499 4320 9563 4324
rect 2044 3836 2108 3840
rect 2044 3780 2048 3836
rect 2048 3780 2104 3836
rect 2104 3780 2108 3836
rect 2044 3776 2108 3780
rect 2124 3836 2188 3840
rect 2124 3780 2128 3836
rect 2128 3780 2184 3836
rect 2184 3780 2188 3836
rect 2124 3776 2188 3780
rect 2204 3836 2268 3840
rect 2204 3780 2208 3836
rect 2208 3780 2264 3836
rect 2264 3780 2268 3836
rect 2204 3776 2268 3780
rect 2284 3836 2348 3840
rect 2284 3780 2288 3836
rect 2288 3780 2344 3836
rect 2344 3780 2348 3836
rect 2284 3776 2348 3780
rect 4229 3836 4293 3840
rect 4229 3780 4233 3836
rect 4233 3780 4289 3836
rect 4289 3780 4293 3836
rect 4229 3776 4293 3780
rect 4309 3836 4373 3840
rect 4309 3780 4313 3836
rect 4313 3780 4369 3836
rect 4369 3780 4373 3836
rect 4309 3776 4373 3780
rect 4389 3836 4453 3840
rect 4389 3780 4393 3836
rect 4393 3780 4449 3836
rect 4449 3780 4453 3836
rect 4389 3776 4453 3780
rect 4469 3836 4533 3840
rect 4469 3780 4473 3836
rect 4473 3780 4529 3836
rect 4529 3780 4533 3836
rect 4469 3776 4533 3780
rect 6414 3836 6478 3840
rect 6414 3780 6418 3836
rect 6418 3780 6474 3836
rect 6474 3780 6478 3836
rect 6414 3776 6478 3780
rect 6494 3836 6558 3840
rect 6494 3780 6498 3836
rect 6498 3780 6554 3836
rect 6554 3780 6558 3836
rect 6494 3776 6558 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 8599 3836 8663 3840
rect 8599 3780 8603 3836
rect 8603 3780 8659 3836
rect 8659 3780 8663 3836
rect 8599 3776 8663 3780
rect 8679 3836 8743 3840
rect 8679 3780 8683 3836
rect 8683 3780 8739 3836
rect 8739 3780 8743 3836
rect 8679 3776 8743 3780
rect 8759 3836 8823 3840
rect 8759 3780 8763 3836
rect 8763 3780 8819 3836
rect 8819 3780 8823 3836
rect 8759 3776 8823 3780
rect 8839 3836 8903 3840
rect 8839 3780 8843 3836
rect 8843 3780 8899 3836
rect 8899 3780 8903 3836
rect 8839 3776 8903 3780
rect 2704 3292 2768 3296
rect 2704 3236 2708 3292
rect 2708 3236 2764 3292
rect 2764 3236 2768 3292
rect 2704 3232 2768 3236
rect 2784 3292 2848 3296
rect 2784 3236 2788 3292
rect 2788 3236 2844 3292
rect 2844 3236 2848 3292
rect 2784 3232 2848 3236
rect 2864 3292 2928 3296
rect 2864 3236 2868 3292
rect 2868 3236 2924 3292
rect 2924 3236 2928 3292
rect 2864 3232 2928 3236
rect 2944 3292 3008 3296
rect 2944 3236 2948 3292
rect 2948 3236 3004 3292
rect 3004 3236 3008 3292
rect 2944 3232 3008 3236
rect 4889 3292 4953 3296
rect 4889 3236 4893 3292
rect 4893 3236 4949 3292
rect 4949 3236 4953 3292
rect 4889 3232 4953 3236
rect 4969 3292 5033 3296
rect 4969 3236 4973 3292
rect 4973 3236 5029 3292
rect 5029 3236 5033 3292
rect 4969 3232 5033 3236
rect 5049 3292 5113 3296
rect 5049 3236 5053 3292
rect 5053 3236 5109 3292
rect 5109 3236 5113 3292
rect 5049 3232 5113 3236
rect 5129 3292 5193 3296
rect 5129 3236 5133 3292
rect 5133 3236 5189 3292
rect 5189 3236 5193 3292
rect 5129 3232 5193 3236
rect 7074 3292 7138 3296
rect 7074 3236 7078 3292
rect 7078 3236 7134 3292
rect 7134 3236 7138 3292
rect 7074 3232 7138 3236
rect 7154 3292 7218 3296
rect 7154 3236 7158 3292
rect 7158 3236 7214 3292
rect 7214 3236 7218 3292
rect 7154 3232 7218 3236
rect 7234 3292 7298 3296
rect 7234 3236 7238 3292
rect 7238 3236 7294 3292
rect 7294 3236 7298 3292
rect 7234 3232 7298 3236
rect 7314 3292 7378 3296
rect 7314 3236 7318 3292
rect 7318 3236 7374 3292
rect 7374 3236 7378 3292
rect 7314 3232 7378 3236
rect 9259 3292 9323 3296
rect 9259 3236 9263 3292
rect 9263 3236 9319 3292
rect 9319 3236 9323 3292
rect 9259 3232 9323 3236
rect 9339 3292 9403 3296
rect 9339 3236 9343 3292
rect 9343 3236 9399 3292
rect 9399 3236 9403 3292
rect 9339 3232 9403 3236
rect 9419 3292 9483 3296
rect 9419 3236 9423 3292
rect 9423 3236 9479 3292
rect 9479 3236 9483 3292
rect 9419 3232 9483 3236
rect 9499 3292 9563 3296
rect 9499 3236 9503 3292
rect 9503 3236 9559 3292
rect 9559 3236 9563 3292
rect 9499 3232 9563 3236
rect 2044 2748 2108 2752
rect 2044 2692 2048 2748
rect 2048 2692 2104 2748
rect 2104 2692 2108 2748
rect 2044 2688 2108 2692
rect 2124 2748 2188 2752
rect 2124 2692 2128 2748
rect 2128 2692 2184 2748
rect 2184 2692 2188 2748
rect 2124 2688 2188 2692
rect 2204 2748 2268 2752
rect 2204 2692 2208 2748
rect 2208 2692 2264 2748
rect 2264 2692 2268 2748
rect 2204 2688 2268 2692
rect 2284 2748 2348 2752
rect 2284 2692 2288 2748
rect 2288 2692 2344 2748
rect 2344 2692 2348 2748
rect 2284 2688 2348 2692
rect 4229 2748 4293 2752
rect 4229 2692 4233 2748
rect 4233 2692 4289 2748
rect 4289 2692 4293 2748
rect 4229 2688 4293 2692
rect 4309 2748 4373 2752
rect 4309 2692 4313 2748
rect 4313 2692 4369 2748
rect 4369 2692 4373 2748
rect 4309 2688 4373 2692
rect 4389 2748 4453 2752
rect 4389 2692 4393 2748
rect 4393 2692 4449 2748
rect 4449 2692 4453 2748
rect 4389 2688 4453 2692
rect 4469 2748 4533 2752
rect 4469 2692 4473 2748
rect 4473 2692 4529 2748
rect 4529 2692 4533 2748
rect 4469 2688 4533 2692
rect 6414 2748 6478 2752
rect 6414 2692 6418 2748
rect 6418 2692 6474 2748
rect 6474 2692 6478 2748
rect 6414 2688 6478 2692
rect 6494 2748 6558 2752
rect 6494 2692 6498 2748
rect 6498 2692 6554 2748
rect 6554 2692 6558 2748
rect 6494 2688 6558 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 8599 2748 8663 2752
rect 8599 2692 8603 2748
rect 8603 2692 8659 2748
rect 8659 2692 8663 2748
rect 8599 2688 8663 2692
rect 8679 2748 8743 2752
rect 8679 2692 8683 2748
rect 8683 2692 8739 2748
rect 8739 2692 8743 2748
rect 8679 2688 8743 2692
rect 8759 2748 8823 2752
rect 8759 2692 8763 2748
rect 8763 2692 8819 2748
rect 8819 2692 8823 2748
rect 8759 2688 8823 2692
rect 8839 2748 8903 2752
rect 8839 2692 8843 2748
rect 8843 2692 8899 2748
rect 8899 2692 8903 2748
rect 8839 2688 8903 2692
rect 2704 2204 2768 2208
rect 2704 2148 2708 2204
rect 2708 2148 2764 2204
rect 2764 2148 2768 2204
rect 2704 2144 2768 2148
rect 2784 2204 2848 2208
rect 2784 2148 2788 2204
rect 2788 2148 2844 2204
rect 2844 2148 2848 2204
rect 2784 2144 2848 2148
rect 2864 2204 2928 2208
rect 2864 2148 2868 2204
rect 2868 2148 2924 2204
rect 2924 2148 2928 2204
rect 2864 2144 2928 2148
rect 2944 2204 3008 2208
rect 2944 2148 2948 2204
rect 2948 2148 3004 2204
rect 3004 2148 3008 2204
rect 2944 2144 3008 2148
rect 4889 2204 4953 2208
rect 4889 2148 4893 2204
rect 4893 2148 4949 2204
rect 4949 2148 4953 2204
rect 4889 2144 4953 2148
rect 4969 2204 5033 2208
rect 4969 2148 4973 2204
rect 4973 2148 5029 2204
rect 5029 2148 5033 2204
rect 4969 2144 5033 2148
rect 5049 2204 5113 2208
rect 5049 2148 5053 2204
rect 5053 2148 5109 2204
rect 5109 2148 5113 2204
rect 5049 2144 5113 2148
rect 5129 2204 5193 2208
rect 5129 2148 5133 2204
rect 5133 2148 5189 2204
rect 5189 2148 5193 2204
rect 5129 2144 5193 2148
rect 7074 2204 7138 2208
rect 7074 2148 7078 2204
rect 7078 2148 7134 2204
rect 7134 2148 7138 2204
rect 7074 2144 7138 2148
rect 7154 2204 7218 2208
rect 7154 2148 7158 2204
rect 7158 2148 7214 2204
rect 7214 2148 7218 2204
rect 7154 2144 7218 2148
rect 7234 2204 7298 2208
rect 7234 2148 7238 2204
rect 7238 2148 7294 2204
rect 7294 2148 7298 2204
rect 7234 2144 7298 2148
rect 7314 2204 7378 2208
rect 7314 2148 7318 2204
rect 7318 2148 7374 2204
rect 7374 2148 7378 2204
rect 7314 2144 7378 2148
rect 9259 2204 9323 2208
rect 9259 2148 9263 2204
rect 9263 2148 9319 2204
rect 9319 2148 9323 2204
rect 9259 2144 9323 2148
rect 9339 2204 9403 2208
rect 9339 2148 9343 2204
rect 9343 2148 9399 2204
rect 9399 2148 9403 2204
rect 9339 2144 9403 2148
rect 9419 2204 9483 2208
rect 9419 2148 9423 2204
rect 9423 2148 9479 2204
rect 9479 2148 9483 2204
rect 9419 2144 9483 2148
rect 9499 2204 9563 2208
rect 9499 2148 9503 2204
rect 9503 2148 9559 2204
rect 9559 2148 9563 2204
rect 9499 2144 9563 2148
<< metal4 >>
rect 2036 10368 2356 10928
rect 2036 10304 2044 10368
rect 2108 10304 2124 10368
rect 2188 10304 2204 10368
rect 2268 10304 2284 10368
rect 2348 10304 2356 10368
rect 2036 9906 2356 10304
rect 2036 9670 2078 9906
rect 2314 9670 2356 9906
rect 2036 9280 2356 9670
rect 2036 9216 2044 9280
rect 2108 9216 2124 9280
rect 2188 9216 2204 9280
rect 2268 9216 2284 9280
rect 2348 9216 2356 9280
rect 2036 8192 2356 9216
rect 2036 8128 2044 8192
rect 2108 8128 2124 8192
rect 2188 8128 2204 8192
rect 2268 8128 2284 8192
rect 2348 8128 2356 8192
rect 2036 7731 2356 8128
rect 2036 7495 2078 7731
rect 2314 7495 2356 7731
rect 2036 7104 2356 7495
rect 2036 7040 2044 7104
rect 2108 7040 2124 7104
rect 2188 7040 2204 7104
rect 2268 7040 2284 7104
rect 2348 7040 2356 7104
rect 2036 6016 2356 7040
rect 2036 5952 2044 6016
rect 2108 5952 2124 6016
rect 2188 5952 2204 6016
rect 2268 5952 2284 6016
rect 2348 5952 2356 6016
rect 2036 5556 2356 5952
rect 2036 5320 2078 5556
rect 2314 5320 2356 5556
rect 2036 4928 2356 5320
rect 2036 4864 2044 4928
rect 2108 4864 2124 4928
rect 2188 4864 2204 4928
rect 2268 4864 2284 4928
rect 2348 4864 2356 4928
rect 2036 3840 2356 4864
rect 2036 3776 2044 3840
rect 2108 3776 2124 3840
rect 2188 3776 2204 3840
rect 2268 3776 2284 3840
rect 2348 3776 2356 3840
rect 2036 3381 2356 3776
rect 2036 3145 2078 3381
rect 2314 3145 2356 3381
rect 2036 2752 2356 3145
rect 2036 2688 2044 2752
rect 2108 2688 2124 2752
rect 2188 2688 2204 2752
rect 2268 2688 2284 2752
rect 2348 2688 2356 2752
rect 2036 2128 2356 2688
rect 2696 10912 3016 10928
rect 2696 10848 2704 10912
rect 2768 10848 2784 10912
rect 2848 10848 2864 10912
rect 2928 10848 2944 10912
rect 3008 10848 3016 10912
rect 2696 10566 3016 10848
rect 2696 10330 2738 10566
rect 2974 10330 3016 10566
rect 2696 9824 3016 10330
rect 2696 9760 2704 9824
rect 2768 9760 2784 9824
rect 2848 9760 2864 9824
rect 2928 9760 2944 9824
rect 3008 9760 3016 9824
rect 2696 8736 3016 9760
rect 2696 8672 2704 8736
rect 2768 8672 2784 8736
rect 2848 8672 2864 8736
rect 2928 8672 2944 8736
rect 3008 8672 3016 8736
rect 2696 8391 3016 8672
rect 2696 8155 2738 8391
rect 2974 8155 3016 8391
rect 2696 7648 3016 8155
rect 2696 7584 2704 7648
rect 2768 7584 2784 7648
rect 2848 7584 2864 7648
rect 2928 7584 2944 7648
rect 3008 7584 3016 7648
rect 2696 6560 3016 7584
rect 2696 6496 2704 6560
rect 2768 6496 2784 6560
rect 2848 6496 2864 6560
rect 2928 6496 2944 6560
rect 3008 6496 3016 6560
rect 2696 6216 3016 6496
rect 2696 5980 2738 6216
rect 2974 5980 3016 6216
rect 2696 5472 3016 5980
rect 2696 5408 2704 5472
rect 2768 5408 2784 5472
rect 2848 5408 2864 5472
rect 2928 5408 2944 5472
rect 3008 5408 3016 5472
rect 2696 4384 3016 5408
rect 2696 4320 2704 4384
rect 2768 4320 2784 4384
rect 2848 4320 2864 4384
rect 2928 4320 2944 4384
rect 3008 4320 3016 4384
rect 2696 4041 3016 4320
rect 2696 3805 2738 4041
rect 2974 3805 3016 4041
rect 2696 3296 3016 3805
rect 2696 3232 2704 3296
rect 2768 3232 2784 3296
rect 2848 3232 2864 3296
rect 2928 3232 2944 3296
rect 3008 3232 3016 3296
rect 2696 2208 3016 3232
rect 2696 2144 2704 2208
rect 2768 2144 2784 2208
rect 2848 2144 2864 2208
rect 2928 2144 2944 2208
rect 3008 2144 3016 2208
rect 2696 2128 3016 2144
rect 4221 10368 4541 10928
rect 4221 10304 4229 10368
rect 4293 10304 4309 10368
rect 4373 10304 4389 10368
rect 4453 10304 4469 10368
rect 4533 10304 4541 10368
rect 4221 9906 4541 10304
rect 4221 9670 4263 9906
rect 4499 9670 4541 9906
rect 4221 9280 4541 9670
rect 4221 9216 4229 9280
rect 4293 9216 4309 9280
rect 4373 9216 4389 9280
rect 4453 9216 4469 9280
rect 4533 9216 4541 9280
rect 4221 8192 4541 9216
rect 4221 8128 4229 8192
rect 4293 8128 4309 8192
rect 4373 8128 4389 8192
rect 4453 8128 4469 8192
rect 4533 8128 4541 8192
rect 4221 7731 4541 8128
rect 4221 7495 4263 7731
rect 4499 7495 4541 7731
rect 4221 7104 4541 7495
rect 4221 7040 4229 7104
rect 4293 7040 4309 7104
rect 4373 7040 4389 7104
rect 4453 7040 4469 7104
rect 4533 7040 4541 7104
rect 4221 6016 4541 7040
rect 4221 5952 4229 6016
rect 4293 5952 4309 6016
rect 4373 5952 4389 6016
rect 4453 5952 4469 6016
rect 4533 5952 4541 6016
rect 4221 5556 4541 5952
rect 4221 5320 4263 5556
rect 4499 5320 4541 5556
rect 4221 4928 4541 5320
rect 4221 4864 4229 4928
rect 4293 4864 4309 4928
rect 4373 4864 4389 4928
rect 4453 4864 4469 4928
rect 4533 4864 4541 4928
rect 4221 3840 4541 4864
rect 4221 3776 4229 3840
rect 4293 3776 4309 3840
rect 4373 3776 4389 3840
rect 4453 3776 4469 3840
rect 4533 3776 4541 3840
rect 4221 3381 4541 3776
rect 4221 3145 4263 3381
rect 4499 3145 4541 3381
rect 4221 2752 4541 3145
rect 4221 2688 4229 2752
rect 4293 2688 4309 2752
rect 4373 2688 4389 2752
rect 4453 2688 4469 2752
rect 4533 2688 4541 2752
rect 4221 2128 4541 2688
rect 4881 10912 5201 10928
rect 4881 10848 4889 10912
rect 4953 10848 4969 10912
rect 5033 10848 5049 10912
rect 5113 10848 5129 10912
rect 5193 10848 5201 10912
rect 4881 10566 5201 10848
rect 4881 10330 4923 10566
rect 5159 10330 5201 10566
rect 4881 9824 5201 10330
rect 4881 9760 4889 9824
rect 4953 9760 4969 9824
rect 5033 9760 5049 9824
rect 5113 9760 5129 9824
rect 5193 9760 5201 9824
rect 4881 8736 5201 9760
rect 4881 8672 4889 8736
rect 4953 8672 4969 8736
rect 5033 8672 5049 8736
rect 5113 8672 5129 8736
rect 5193 8672 5201 8736
rect 4881 8391 5201 8672
rect 4881 8155 4923 8391
rect 5159 8155 5201 8391
rect 4881 7648 5201 8155
rect 4881 7584 4889 7648
rect 4953 7584 4969 7648
rect 5033 7584 5049 7648
rect 5113 7584 5129 7648
rect 5193 7584 5201 7648
rect 4881 6560 5201 7584
rect 4881 6496 4889 6560
rect 4953 6496 4969 6560
rect 5033 6496 5049 6560
rect 5113 6496 5129 6560
rect 5193 6496 5201 6560
rect 4881 6216 5201 6496
rect 4881 5980 4923 6216
rect 5159 5980 5201 6216
rect 4881 5472 5201 5980
rect 4881 5408 4889 5472
rect 4953 5408 4969 5472
rect 5033 5408 5049 5472
rect 5113 5408 5129 5472
rect 5193 5408 5201 5472
rect 4881 4384 5201 5408
rect 4881 4320 4889 4384
rect 4953 4320 4969 4384
rect 5033 4320 5049 4384
rect 5113 4320 5129 4384
rect 5193 4320 5201 4384
rect 4881 4041 5201 4320
rect 4881 3805 4923 4041
rect 5159 3805 5201 4041
rect 4881 3296 5201 3805
rect 4881 3232 4889 3296
rect 4953 3232 4969 3296
rect 5033 3232 5049 3296
rect 5113 3232 5129 3296
rect 5193 3232 5201 3296
rect 4881 2208 5201 3232
rect 4881 2144 4889 2208
rect 4953 2144 4969 2208
rect 5033 2144 5049 2208
rect 5113 2144 5129 2208
rect 5193 2144 5201 2208
rect 4881 2128 5201 2144
rect 6406 10368 6726 10928
rect 6406 10304 6414 10368
rect 6478 10304 6494 10368
rect 6558 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6726 10368
rect 6406 9906 6726 10304
rect 6406 9670 6448 9906
rect 6684 9670 6726 9906
rect 6406 9280 6726 9670
rect 6406 9216 6414 9280
rect 6478 9216 6494 9280
rect 6558 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6726 9280
rect 6406 8192 6726 9216
rect 6406 8128 6414 8192
rect 6478 8128 6494 8192
rect 6558 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6726 8192
rect 6406 7731 6726 8128
rect 6406 7495 6448 7731
rect 6684 7495 6726 7731
rect 6406 7104 6726 7495
rect 6406 7040 6414 7104
rect 6478 7040 6494 7104
rect 6558 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6726 7104
rect 6406 6016 6726 7040
rect 6406 5952 6414 6016
rect 6478 5952 6494 6016
rect 6558 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6726 6016
rect 6406 5556 6726 5952
rect 6406 5320 6448 5556
rect 6684 5320 6726 5556
rect 6406 4928 6726 5320
rect 6406 4864 6414 4928
rect 6478 4864 6494 4928
rect 6558 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6726 4928
rect 6406 3840 6726 4864
rect 6406 3776 6414 3840
rect 6478 3776 6494 3840
rect 6558 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6726 3840
rect 6406 3381 6726 3776
rect 6406 3145 6448 3381
rect 6684 3145 6726 3381
rect 6406 2752 6726 3145
rect 6406 2688 6414 2752
rect 6478 2688 6494 2752
rect 6558 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6726 2752
rect 6406 2128 6726 2688
rect 7066 10912 7386 10928
rect 7066 10848 7074 10912
rect 7138 10848 7154 10912
rect 7218 10848 7234 10912
rect 7298 10848 7314 10912
rect 7378 10848 7386 10912
rect 7066 10566 7386 10848
rect 7066 10330 7108 10566
rect 7344 10330 7386 10566
rect 7066 9824 7386 10330
rect 7066 9760 7074 9824
rect 7138 9760 7154 9824
rect 7218 9760 7234 9824
rect 7298 9760 7314 9824
rect 7378 9760 7386 9824
rect 7066 8736 7386 9760
rect 7066 8672 7074 8736
rect 7138 8672 7154 8736
rect 7218 8672 7234 8736
rect 7298 8672 7314 8736
rect 7378 8672 7386 8736
rect 7066 8391 7386 8672
rect 7066 8155 7108 8391
rect 7344 8155 7386 8391
rect 7066 7648 7386 8155
rect 7066 7584 7074 7648
rect 7138 7584 7154 7648
rect 7218 7584 7234 7648
rect 7298 7584 7314 7648
rect 7378 7584 7386 7648
rect 7066 6560 7386 7584
rect 7066 6496 7074 6560
rect 7138 6496 7154 6560
rect 7218 6496 7234 6560
rect 7298 6496 7314 6560
rect 7378 6496 7386 6560
rect 7066 6216 7386 6496
rect 7066 5980 7108 6216
rect 7344 5980 7386 6216
rect 7066 5472 7386 5980
rect 7066 5408 7074 5472
rect 7138 5408 7154 5472
rect 7218 5408 7234 5472
rect 7298 5408 7314 5472
rect 7378 5408 7386 5472
rect 7066 4384 7386 5408
rect 7066 4320 7074 4384
rect 7138 4320 7154 4384
rect 7218 4320 7234 4384
rect 7298 4320 7314 4384
rect 7378 4320 7386 4384
rect 7066 4041 7386 4320
rect 7066 3805 7108 4041
rect 7344 3805 7386 4041
rect 7066 3296 7386 3805
rect 7066 3232 7074 3296
rect 7138 3232 7154 3296
rect 7218 3232 7234 3296
rect 7298 3232 7314 3296
rect 7378 3232 7386 3296
rect 7066 2208 7386 3232
rect 7066 2144 7074 2208
rect 7138 2144 7154 2208
rect 7218 2144 7234 2208
rect 7298 2144 7314 2208
rect 7378 2144 7386 2208
rect 7066 2128 7386 2144
rect 8591 10368 8911 10928
rect 8591 10304 8599 10368
rect 8663 10304 8679 10368
rect 8743 10304 8759 10368
rect 8823 10304 8839 10368
rect 8903 10304 8911 10368
rect 8591 9906 8911 10304
rect 8591 9670 8633 9906
rect 8869 9670 8911 9906
rect 8591 9280 8911 9670
rect 8591 9216 8599 9280
rect 8663 9216 8679 9280
rect 8743 9216 8759 9280
rect 8823 9216 8839 9280
rect 8903 9216 8911 9280
rect 8591 8192 8911 9216
rect 8591 8128 8599 8192
rect 8663 8128 8679 8192
rect 8743 8128 8759 8192
rect 8823 8128 8839 8192
rect 8903 8128 8911 8192
rect 8591 7731 8911 8128
rect 8591 7495 8633 7731
rect 8869 7495 8911 7731
rect 8591 7104 8911 7495
rect 8591 7040 8599 7104
rect 8663 7040 8679 7104
rect 8743 7040 8759 7104
rect 8823 7040 8839 7104
rect 8903 7040 8911 7104
rect 8591 6016 8911 7040
rect 8591 5952 8599 6016
rect 8663 5952 8679 6016
rect 8743 5952 8759 6016
rect 8823 5952 8839 6016
rect 8903 5952 8911 6016
rect 8591 5556 8911 5952
rect 8591 5320 8633 5556
rect 8869 5320 8911 5556
rect 8591 4928 8911 5320
rect 8591 4864 8599 4928
rect 8663 4864 8679 4928
rect 8743 4864 8759 4928
rect 8823 4864 8839 4928
rect 8903 4864 8911 4928
rect 8591 3840 8911 4864
rect 8591 3776 8599 3840
rect 8663 3776 8679 3840
rect 8743 3776 8759 3840
rect 8823 3776 8839 3840
rect 8903 3776 8911 3840
rect 8591 3381 8911 3776
rect 8591 3145 8633 3381
rect 8869 3145 8911 3381
rect 8591 2752 8911 3145
rect 8591 2688 8599 2752
rect 8663 2688 8679 2752
rect 8743 2688 8759 2752
rect 8823 2688 8839 2752
rect 8903 2688 8911 2752
rect 8591 2128 8911 2688
rect 9251 10912 9571 10928
rect 9251 10848 9259 10912
rect 9323 10848 9339 10912
rect 9403 10848 9419 10912
rect 9483 10848 9499 10912
rect 9563 10848 9571 10912
rect 9251 10566 9571 10848
rect 9251 10330 9293 10566
rect 9529 10330 9571 10566
rect 9251 9824 9571 10330
rect 9251 9760 9259 9824
rect 9323 9760 9339 9824
rect 9403 9760 9419 9824
rect 9483 9760 9499 9824
rect 9563 9760 9571 9824
rect 9251 8736 9571 9760
rect 9251 8672 9259 8736
rect 9323 8672 9339 8736
rect 9403 8672 9419 8736
rect 9483 8672 9499 8736
rect 9563 8672 9571 8736
rect 9251 8391 9571 8672
rect 9251 8155 9293 8391
rect 9529 8155 9571 8391
rect 9251 7648 9571 8155
rect 9251 7584 9259 7648
rect 9323 7584 9339 7648
rect 9403 7584 9419 7648
rect 9483 7584 9499 7648
rect 9563 7584 9571 7648
rect 9251 6560 9571 7584
rect 9251 6496 9259 6560
rect 9323 6496 9339 6560
rect 9403 6496 9419 6560
rect 9483 6496 9499 6560
rect 9563 6496 9571 6560
rect 9251 6216 9571 6496
rect 9251 5980 9293 6216
rect 9529 5980 9571 6216
rect 9251 5472 9571 5980
rect 9251 5408 9259 5472
rect 9323 5408 9339 5472
rect 9403 5408 9419 5472
rect 9483 5408 9499 5472
rect 9563 5408 9571 5472
rect 9251 4384 9571 5408
rect 9251 4320 9259 4384
rect 9323 4320 9339 4384
rect 9403 4320 9419 4384
rect 9483 4320 9499 4384
rect 9563 4320 9571 4384
rect 9251 4041 9571 4320
rect 9251 3805 9293 4041
rect 9529 3805 9571 4041
rect 9251 3296 9571 3805
rect 9251 3232 9259 3296
rect 9323 3232 9339 3296
rect 9403 3232 9419 3296
rect 9483 3232 9499 3296
rect 9563 3232 9571 3296
rect 9251 2208 9571 3232
rect 9251 2144 9259 2208
rect 9323 2144 9339 2208
rect 9403 2144 9419 2208
rect 9483 2144 9499 2208
rect 9563 2144 9571 2208
rect 9251 2128 9571 2144
<< via4 >>
rect 2078 9670 2314 9906
rect 2078 7495 2314 7731
rect 2078 5320 2314 5556
rect 2078 3145 2314 3381
rect 2738 10330 2974 10566
rect 2738 8155 2974 8391
rect 2738 5980 2974 6216
rect 2738 3805 2974 4041
rect 4263 9670 4499 9906
rect 4263 7495 4499 7731
rect 4263 5320 4499 5556
rect 4263 3145 4499 3381
rect 4923 10330 5159 10566
rect 4923 8155 5159 8391
rect 4923 5980 5159 6216
rect 4923 3805 5159 4041
rect 6448 9670 6684 9906
rect 6448 7495 6684 7731
rect 6448 5320 6684 5556
rect 6448 3145 6684 3381
rect 7108 10330 7344 10566
rect 7108 8155 7344 8391
rect 7108 5980 7344 6216
rect 7108 3805 7344 4041
rect 8633 9670 8869 9906
rect 8633 7495 8869 7731
rect 8633 5320 8869 5556
rect 8633 3145 8869 3381
rect 9293 10330 9529 10566
rect 9293 8155 9529 8391
rect 9293 5980 9529 6216
rect 9293 3805 9529 4041
<< metal5 >>
rect 1056 10566 9892 10608
rect 1056 10330 2738 10566
rect 2974 10330 4923 10566
rect 5159 10330 7108 10566
rect 7344 10330 9293 10566
rect 9529 10330 9892 10566
rect 1056 10288 9892 10330
rect 1056 9906 9892 9948
rect 1056 9670 2078 9906
rect 2314 9670 4263 9906
rect 4499 9670 6448 9906
rect 6684 9670 8633 9906
rect 8869 9670 9892 9906
rect 1056 9628 9892 9670
rect 1056 8391 9892 8433
rect 1056 8155 2738 8391
rect 2974 8155 4923 8391
rect 5159 8155 7108 8391
rect 7344 8155 9293 8391
rect 9529 8155 9892 8391
rect 1056 8113 9892 8155
rect 1056 7731 9892 7773
rect 1056 7495 2078 7731
rect 2314 7495 4263 7731
rect 4499 7495 6448 7731
rect 6684 7495 8633 7731
rect 8869 7495 9892 7731
rect 1056 7453 9892 7495
rect 1056 6216 9892 6258
rect 1056 5980 2738 6216
rect 2974 5980 4923 6216
rect 5159 5980 7108 6216
rect 7344 5980 9293 6216
rect 9529 5980 9892 6216
rect 1056 5938 9892 5980
rect 1056 5556 9892 5598
rect 1056 5320 2078 5556
rect 2314 5320 4263 5556
rect 4499 5320 6448 5556
rect 6684 5320 8633 5556
rect 8869 5320 9892 5556
rect 1056 5278 9892 5320
rect 1056 4041 9892 4083
rect 1056 3805 2738 4041
rect 2974 3805 4923 4041
rect 5159 3805 7108 4041
rect 7344 3805 9293 4041
rect 9529 3805 9892 4041
rect 1056 3763 9892 3805
rect 1056 3381 9892 3423
rect 1056 3145 2078 3381
rect 2314 3145 4263 3381
rect 4499 3145 6448 3381
rect 6684 3145 8633 3381
rect 8869 3145 9892 3381
rect 1056 3103 9892 3145
use sky130_fd_sc_hd__nor2_4  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7544 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _114_
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_4  _115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__xnor2_4  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 -1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 1704896540
transform -1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 1704896540
transform -1 0 7360 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _120_
timestamp 1704896540
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _121_
timestamp 1704896540
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _123_
timestamp 1704896540
transform 1 0 6900 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6164 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6164 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _130_
timestamp 1704896540
transform 1 0 7544 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _132_
timestamp 1704896540
transform -1 0 8740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _133_
timestamp 1704896540
transform -1 0 8740 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _134_
timestamp 1704896540
transform -1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _137_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1704896540
transform -1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _140_
timestamp 1704896540
transform 1 0 8004 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 1704896540
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _143_
timestamp 1704896540
transform 1 0 8372 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1704896540
transform -1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _145_
timestamp 1704896540
transform 1 0 7636 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7084 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_2  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6164 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _148_
timestamp 1704896540
transform -1 0 5980 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _149_
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _150_
timestamp 1704896540
transform 1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _151_
timestamp 1704896540
transform -1 0 6256 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _152_
timestamp 1704896540
transform -1 0 5888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _153_
timestamp 1704896540
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _154_
timestamp 1704896540
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _155_
timestamp 1704896540
transform -1 0 6808 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _157_
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _158_
timestamp 1704896540
transform -1 0 5520 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3680 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _160_
timestamp 1704896540
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2852 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _163_
timestamp 1704896540
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _164_
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _165_
timestamp 1704896540
transform 1 0 2208 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _166_
timestamp 1704896540
transform -1 0 2208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _167_
timestamp 1704896540
transform -1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1704896540
transform 1 0 3772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4416 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1704896540
transform -1 0 5152 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1704896540
transform 1 0 4048 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 1704896540
transform -1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _176_
timestamp 1704896540
transform -1 0 2576 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _177_
timestamp 1704896540
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _178_
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _179_
timestamp 1704896540
transform -1 0 3496 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _180_
timestamp 1704896540
transform 1 0 2024 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _181_
timestamp 1704896540
transform -1 0 2024 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _182_
timestamp 1704896540
transform -1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1704896540
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _184_
timestamp 1704896540
transform 1 0 4232 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _185_
timestamp 1704896540
transform 1 0 3036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _186_
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _187_
timestamp 1704896540
transform -1 0 3036 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _188_
timestamp 1704896540
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _189_
timestamp 1704896540
transform -1 0 2576 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _190_
timestamp 1704896540
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 1704896540
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _192_
timestamp 1704896540
transform -1 0 3312 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _193_
timestamp 1704896540
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _194_
timestamp 1704896540
transform -1 0 2208 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _195_
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1704896540
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _197_
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _198_
timestamp 1704896540
transform -1 0 3680 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _199_
timestamp 1704896540
transform 1 0 3128 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_4  _200_
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _201_
timestamp 1704896540
transform 1 0 4508 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _202_
timestamp 1704896540
transform -1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _204_
timestamp 1704896540
transform 1 0 4600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _205_
timestamp 1704896540
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _206_
timestamp 1704896540
transform 1 0 4968 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _207_
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _209_
timestamp 1704896540
transform 1 0 5428 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _210_
timestamp 1704896540
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1704896540
transform 1 0 4508 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _214_
timestamp 1704896540
transform 1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _215_
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _216_
timestamp 1704896540
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1704896540
transform -1 0 7268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1704896540
transform 1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1704896540
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1704896540
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1704896540
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1704896540
transform -1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_79
timestamp 1704896540
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_91
timestamp 1704896540
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_21
timestamp 1704896540
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_25
timestamp 1704896540
transform 1 0 3404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_65
timestamp 1704896540
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_84
timestamp 1704896540
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_91
timestamp 1704896540
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_35
timestamp 1704896540
transform 1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 1704896540
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_55
timestamp 1704896540
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_59
timestamp 1704896540
transform 1 0 6532 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 1704896540
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_18
timestamp 1704896540
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_30
timestamp 1704896540
transform 1 0 3864 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_45
timestamp 1704896540
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_66
timestamp 1704896540
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_91
timestamp 1704896540
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_12
timestamp 1704896540
transform 1 0 2208 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_18
timestamp 1704896540
transform 1 0 2760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_38
timestamp 1704896540
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_45
timestamp 1704896540
transform 1 0 5244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_57
timestamp 1704896540
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_19
timestamp 1704896540
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_35
timestamp 1704896540
transform 1 0 4324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_62
timestamp 1704896540
transform 1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_9
timestamp 1704896540
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_21
timestamp 1704896540
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_33
timestamp 1704896540
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_68
timestamp 1704896540
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_90
timestamp 1704896540
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_14
timestamp 1704896540
transform 1 0 2392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_22
timestamp 1704896540
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_36
timestamp 1704896540
transform 1 0 4416 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_78
timestamp 1704896540
transform 1 0 8280 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_39
timestamp 1704896540
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_48
timestamp 1704896540
transform 1 0 5520 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_60
timestamp 1704896540
transform 1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_66
timestamp 1704896540
transform 1 0 7176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_78
timestamp 1704896540
transform 1 0 8280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_10
timestamp 1704896540
transform 1 0 2024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_16
timestamp 1704896540
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_20
timestamp 1704896540
transform 1 0 2944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_37
timestamp 1704896540
transform 1 0 4508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_41
timestamp 1704896540
transform 1 0 4876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_50
timestamp 1704896540
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_67
timestamp 1704896540
transform 1 0 7268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_75
timestamp 1704896540
transform 1 0 8004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 1704896540
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1704896540
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1704896540
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_37
timestamp 1704896540
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_52
timestamp 1704896540
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_20
timestamp 1704896540
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_28
timestamp 1704896540
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_38
timestamp 1704896540
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_42
timestamp 1704896540
transform 1 0 4968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1704896540
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_62
timestamp 1704896540
transform 1 0 6808 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_68
timestamp 1704896540
transform 1 0 7360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_18
timestamp 1704896540
transform 1 0 2760 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_24
timestamp 1704896540
transform 1 0 3312 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_34
timestamp 1704896540
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_42
timestamp 1704896540
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_56
timestamp 1704896540
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_68
timestamp 1704896540
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_74
timestamp 1704896540
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1704896540
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_91
timestamp 1704896540
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_11
timestamp 1704896540
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_23
timestamp 1704896540
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_28
timestamp 1704896540
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_67
timestamp 1704896540
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_6
timestamp 1704896540
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_18
timestamp 1704896540
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_62
timestamp 1704896540
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_79
timestamp 1704896540
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_88
timestamp 1704896540
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_15
timestamp 1704896540
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_66
timestamp 1704896540
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_70
timestamp 1704896540
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_83
timestamp 1704896540
transform 1 0 8740 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_91
timestamp 1704896540
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 9476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 4416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1704896540
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1704896540
transform -1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1704896540
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1704896540
transform -1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1704896540
transform -1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input20
timestamp 1704896540
transform -1 0 9568 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output21
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1704896540
transform -1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1704896540
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1704896540
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output29
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_16
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_17
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_18
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_19
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_20
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_21
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_22
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_23
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_24
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_25
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_26
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_27
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_28
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_29
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_30
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_31
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4968 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 1704896540
transform 1 0 5336 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer4
timestamp 1704896540
transform 1 0 5336 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer5
timestamp 1704896540
transform 1 0 8280 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer6
timestamp 1704896540
transform -1 0 8280 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 1704896540
transform -1 0 4692 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer8
timestamp 1704896540
transform -1 0 8280 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 1704896540
transform -1 0 8280 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer10
timestamp 1704896540
transform 1 0 8096 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer11
timestamp 1704896540
transform -1 0 8832 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer12
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer13
timestamp 1704896540
transform -1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer14
timestamp 1704896540
transform -1 0 3680 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer15
timestamp 1704896540
transform -1 0 5520 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer16
timestamp 1704896540
transform -1 0 5336 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer17
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_35
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_38
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_39
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_40
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_41
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_42
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_43
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_44
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_45
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_46
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_47
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_48
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_49
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_50
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_51
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_52
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_53
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_54
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_55
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_56
timestamp 1704896540
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_57
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1704896540
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 2696 2128 3016 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4881 2128 5201 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7066 2128 7386 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9251 2128 9571 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3763 9892 4083 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5938 9892 6258 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8113 9892 8433 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10288 9892 10608 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2036 2128 2356 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4221 2128 4541 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6406 2128 6726 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8591 2128 8911 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3103 9892 3423 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5278 9892 5598 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7453 9892 7773 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 9628 9892 9948 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 a[0]
port 2 nsew signal input
flabel metal3 s 10164 4768 10964 4888 0 FreeSans 480 0 0 0 a[1]
port 3 nsew signal input
flabel metal2 s 7746 12308 7802 13108 0 FreeSans 224 90 0 0 a[2]
port 4 nsew signal input
flabel metal2 s 6458 12308 6514 13108 0 FreeSans 224 90 0 0 a[3]
port 5 nsew signal input
flabel metal2 s 3882 12308 3938 13108 0 FreeSans 224 90 0 0 a[4]
port 6 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 a[5]
port 7 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 a[6]
port 8 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 a[7]
port 9 nsew signal input
flabel metal3 s 10164 4088 10964 4208 0 FreeSans 480 0 0 0 b[0]
port 10 nsew signal input
flabel metal3 s 10164 5448 10964 5568 0 FreeSans 480 0 0 0 b[1]
port 11 nsew signal input
flabel metal2 s 8390 12308 8446 13108 0 FreeSans 224 90 0 0 b[2]
port 12 nsew signal input
flabel metal2 s 5814 12308 5870 13108 0 FreeSans 224 90 0 0 b[3]
port 13 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 b[4]
port 14 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 b[5]
port 15 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 b[6]
port 16 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 b[7]
port 17 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 cin
port 18 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 cout
port 19 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 op[0]
port 20 nsew signal input
flabel metal3 s 10164 6808 10964 6928 0 FreeSans 480 0 0 0 op[1]
port 21 nsew signal input
flabel metal3 s 10164 8168 10964 8288 0 FreeSans 480 0 0 0 op[2]
port 22 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 result[0]
port 23 nsew signal output
flabel metal3 s 10164 6128 10964 6248 0 FreeSans 480 0 0 0 result[1]
port 24 nsew signal output
flabel metal3 s 10164 7488 10964 7608 0 FreeSans 480 0 0 0 result[2]
port 25 nsew signal output
flabel metal2 s 5170 12308 5226 13108 0 FreeSans 224 90 0 0 result[3]
port 26 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 result[4]
port 27 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 result[5]
port 28 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 result[6]
port 29 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 result[7]
port 30 nsew signal output
rlabel metal1 5474 10880 5474 10880 0 VGND
rlabel metal1 5474 10336 5474 10336 0 VPWR
rlabel metal1 2645 7378 2645 7378 0 _000_
rlabel metal1 2024 6358 2024 6358 0 _001_
rlabel metal2 2162 6460 2162 6460 0 _002_
rlabel metal1 3601 7514 3601 7514 0 _003_
rlabel metal1 3358 6630 3358 6630 0 _004_
rlabel via1 1873 6358 1873 6358 0 _005_
rlabel metal2 1702 6460 1702 6460 0 _006_
rlabel metal1 4554 5712 4554 5712 0 _007_
rlabel metal2 3358 5270 3358 5270 0 _008_
rlabel metal2 4186 6647 4186 6647 0 _009_
rlabel metal2 2622 3162 2622 3162 0 _010_
rlabel metal1 2622 3604 2622 3604 0 _011_
rlabel metal1 2530 3570 2530 3570 0 _012_
rlabel metal1 2070 3366 2070 3366 0 _013_
rlabel metal1 1748 3706 1748 3706 0 _014_
rlabel metal2 2438 4862 2438 4862 0 _015_
rlabel metal1 2852 4794 2852 4794 0 _016_
rlabel metal1 2047 5270 2047 5270 0 _017_
rlabel metal1 1840 4794 1840 4794 0 _018_
rlabel metal2 3266 3332 3266 3332 0 _019_
rlabel metal1 3634 3502 3634 3502 0 _020_
rlabel metal1 4186 3706 4186 3706 0 _021_
rlabel metal1 4186 4590 4186 4590 0 _022_
rlabel metal1 4600 3434 4600 3434 0 _023_
rlabel metal1 5198 3162 5198 3162 0 _024_
rlabel metal1 4324 2822 4324 2822 0 _025_
rlabel metal1 5796 3094 5796 3094 0 _026_
rlabel metal1 5244 3978 5244 3978 0 _027_
rlabel metal1 5014 3910 5014 3910 0 _028_
rlabel metal2 5382 4420 5382 4420 0 _029_
rlabel metal2 5014 4794 5014 4794 0 _030_
rlabel metal1 5566 4794 5566 4794 0 _031_
rlabel metal1 6348 2958 6348 2958 0 _032_
rlabel metal1 5842 3604 5842 3604 0 _033_
rlabel metal1 6578 3162 6578 3162 0 _034_
rlabel metal1 6946 3536 6946 3536 0 _035_
rlabel metal1 6762 4046 6762 4046 0 _036_
rlabel metal1 6946 4114 6946 4114 0 _037_
rlabel metal1 6486 3706 6486 3706 0 _038_
rlabel metal1 1978 6256 1978 6256 0 _039_
rlabel metal1 7590 2992 7590 2992 0 _040_
rlabel metal1 7728 3026 7728 3026 0 _041_
rlabel metal1 7314 3468 7314 3468 0 _042_
rlabel metal2 6210 3264 6210 3264 0 _043_
rlabel metal2 7866 3332 7866 3332 0 _044_
rlabel metal1 8556 3162 8556 3162 0 _045_
rlabel metal2 6394 5338 6394 5338 0 _046_
rlabel metal1 9430 6698 9430 6698 0 _047_
rlabel metal1 9614 3570 9614 3570 0 _048_
rlabel metal2 8418 4386 8418 4386 0 _049_
rlabel metal2 8234 5372 8234 5372 0 _050_
rlabel metal1 7130 5338 7130 5338 0 _051_
rlabel metal1 5934 5712 5934 5712 0 _052_
rlabel metal1 1564 6698 1564 6698 0 _053_
rlabel metal2 6762 4590 6762 4590 0 _054_
rlabel metal1 6026 5338 6026 5338 0 _055_
rlabel metal1 8096 5882 8096 5882 0 _056_
rlabel metal1 8602 7888 8602 7888 0 _057_
rlabel metal1 6578 7854 6578 7854 0 _058_
rlabel metal2 2622 7582 2622 7582 0 _059_
rlabel metal1 5474 5780 5474 5780 0 _060_
rlabel metal2 8510 5372 8510 5372 0 _061_
rlabel metal1 8234 7310 8234 7310 0 _062_
rlabel metal1 7958 5814 7958 5814 0 _063_
rlabel metal1 9016 7854 9016 7854 0 _064_
rlabel metal1 8648 9894 8648 9894 0 _065_
rlabel metal2 8326 10049 8326 10049 0 _066_
rlabel metal1 9522 9350 9522 9350 0 _067_
rlabel metal1 8418 8262 8418 8262 0 _068_
rlabel metal2 8970 7888 8970 7888 0 _069_
rlabel metal1 8050 7922 8050 7922 0 _070_
rlabel metal1 7912 7990 7912 7990 0 _071_
rlabel metal2 8510 8636 8510 8636 0 _072_
rlabel metal1 8004 8058 8004 8058 0 _073_
rlabel metal1 9016 9486 9016 9486 0 _074_
rlabel metal2 8418 9826 8418 9826 0 _075_
rlabel via1 8155 9622 8155 9622 0 _076_
rlabel metal1 7728 9690 7728 9690 0 _077_
rlabel metal1 6348 9962 6348 9962 0 _078_
rlabel metal1 5244 10098 5244 10098 0 _079_
rlabel metal1 5290 7344 5290 7344 0 _080_
rlabel metal1 5198 7412 5198 7412 0 _081_
rlabel metal1 6762 8432 6762 8432 0 _082_
rlabel metal2 5474 8908 5474 8908 0 _083_
rlabel metal1 5681 7446 5681 7446 0 _084_
rlabel metal2 5658 7820 5658 7820 0 _085_
rlabel metal1 6026 9622 6026 9622 0 _086_
rlabel metal1 3496 9690 3496 9690 0 _087_
rlabel metal1 5290 8500 5290 8500 0 _088_
rlabel metal1 4876 8942 4876 8942 0 _089_
rlabel metal1 3542 10642 3542 10642 0 _090_
rlabel metal1 3220 9350 3220 9350 0 _091_
rlabel metal1 2162 8976 2162 8976 0 _092_
rlabel metal1 2254 8908 2254 8908 0 _093_
rlabel metal2 2530 8772 2530 8772 0 _094_
rlabel metal2 3818 8636 3818 8636 0 _095_
rlabel metal1 2116 8602 2116 8602 0 _096_
rlabel metal2 1794 8772 1794 8772 0 _097_
rlabel metal1 4002 9554 4002 9554 0 _098_
rlabel metal1 4554 9146 4554 9146 0 _099_
rlabel metal2 4278 7565 4278 7565 0 _100_
rlabel metal1 4554 8466 4554 8466 0 _101_
rlabel metal1 4148 7514 4148 7514 0 _102_
rlabel metal1 4738 5712 4738 5712 0 _103_
rlabel metal1 4462 5644 4462 5644 0 _104_
rlabel metal2 8418 1588 8418 1588 0 a[0]
rlabel metal1 9522 4114 9522 4114 0 a[1]
rlabel metal1 9430 10676 9430 10676 0 a[2]
rlabel metal1 6762 10642 6762 10642 0 a[3]
rlabel metal1 4462 10676 4462 10676 0 a[4]
rlabel metal3 751 7548 751 7548 0 a[5]
rlabel metal2 3266 1588 3266 1588 0 a[6]
rlabel metal2 3910 1588 3910 1588 0 a[7]
rlabel metal1 7314 3366 7314 3366 0 alu0.result
rlabel metal2 6118 6086 6118 6086 0 alu1.result
rlabel metal1 8832 8058 8832 8058 0 alu2.result
rlabel metal1 4830 7514 4830 7514 0 alu3.result
rlabel metal1 2576 8942 2576 8942 0 alu4.result
rlabel metal1 2392 6426 2392 6426 0 alu5.result
rlabel metal1 1472 5338 1472 5338 0 alu6.result
rlabel metal1 4600 5202 4600 5202 0 alu7.result
rlabel metal1 6578 4624 6578 4624 0 b[0]
rlabel via2 7222 5219 7222 5219 0 b[1]
rlabel metal1 8970 10064 8970 10064 0 b[2]
rlabel metal1 5934 10642 5934 10642 0 b[3]
rlabel metal3 1050 9588 1050 9588 0 b[4]
rlabel metal3 1050 5508 1050 5508 0 b[5]
rlabel metal3 1050 4148 1050 4148 0 b[6]
rlabel metal2 5198 1027 5198 1027 0 b[7]
rlabel metal2 7774 1520 7774 1520 0 cin
rlabel metal2 5842 1554 5842 1554 0 cout
rlabel metal1 7590 4556 7590 4556 0 net1
rlabel metal1 7130 5712 7130 5712 0 net10
rlabel metal1 8924 10642 8924 10642 0 net11
rlabel metal1 5750 8432 5750 8432 0 net12
rlabel metal2 2622 9724 2622 9724 0 net13
rlabel metal1 2806 6834 2806 6834 0 net14
rlabel metal1 2116 3570 2116 3570 0 net15
rlabel metal1 5382 2618 5382 2618 0 net16
rlabel metal1 8050 2448 8050 2448 0 net17
rlabel metal1 5014 6222 5014 6222 0 net18
rlabel metal1 8234 7378 8234 7378 0 net19
rlabel metal1 8740 3910 8740 3910 0 net2
rlabel metal2 8418 8738 8418 8738 0 net20
rlabel metal1 6394 2414 6394 2414 0 net21
rlabel metal1 7544 2414 7544 2414 0 net22
rlabel metal1 7268 6290 7268 6290 0 net23
rlabel metal2 7590 7922 7590 7922 0 net24
rlabel metal1 5474 8058 5474 8058 0 net25
rlabel metal1 1702 8874 1702 8874 0 net26
rlabel metal1 1748 7378 1748 7378 0 net27
rlabel metal2 1702 5066 1702 5066 0 net28
rlabel metal2 4738 3757 4738 3757 0 net29
rlabel metal1 8418 9554 8418 9554 0 net3
rlabel metal1 4186 10098 4186 10098 0 net30
rlabel metal1 3634 9520 3634 9520 0 net31
rlabel metal1 5612 9010 5612 9010 0 net32
rlabel metal1 4922 7888 4922 7888 0 net33
rlabel metal2 8142 4930 8142 4930 0 net34
rlabel metal1 4968 6766 4968 6766 0 net35
rlabel metal1 4462 4658 4462 4658 0 net36
rlabel metal1 8004 10098 8004 10098 0 net37
rlabel metal2 6946 10030 6946 10030 0 net38
rlabel metal2 9246 7004 9246 7004 0 net39
rlabel metal1 6808 10030 6808 10030 0 net4
rlabel metal1 7820 5610 7820 5610 0 net40
rlabel metal2 9154 7276 9154 7276 0 net41
rlabel metal1 5934 3672 5934 3672 0 net42
rlabel metal2 3174 9724 3174 9724 0 net43
rlabel metal1 7590 10132 7590 10132 0 net44
rlabel metal1 3910 10608 3910 10608 0 net45
rlabel metal1 6854 6188 6854 6188 0 net46
rlabel metal1 3634 8908 3634 8908 0 net5
rlabel metal2 3818 7548 3818 7548 0 net6
rlabel metal1 3174 2618 3174 2618 0 net7
rlabel metal1 4646 3026 4646 3026 0 net8
rlabel metal1 7360 3026 7360 3026 0 net9
rlabel metal3 751 6188 751 6188 0 op[0]
rlabel metal2 9430 7123 9430 7123 0 op[1]
rlabel metal2 9430 8347 9430 8347 0 op[2]
rlabel metal2 7130 959 7130 959 0 result[0]
rlabel via2 7498 6171 7498 6171 0 result[1]
rlabel metal2 7406 7021 7406 7021 0 result[2]
rlabel metal1 5934 10778 5934 10778 0 result[3]
rlabel metal3 751 8908 751 8908 0 result[4]
rlabel metal3 1096 6868 1096 6868 0 result[5]
rlabel metal1 1380 4794 1380 4794 0 result[6]
rlabel metal2 4554 1554 4554 1554 0 result[7]
<< properties >>
string FIXED_BBOX 0 0 10964 13108
<< end >>
